magic
tech sky130B
magscale 1 2
timestamp 1675206000
<< checkpaint >>
rect 0 0 50448 15816
<< m2 >>
rect 0 924 48600 1076
rect 924 924 49524 1076
rect 0 12740 48600 12892
rect 924 12740 49524 12892
rect 1384 13768 34632 13920
rect 1384 13768 34632 13920
rect 9160 14208 26856 14360
rect 9160 14208 26856 14360
rect 40264 14432 40464 14584
rect 40264 14432 40464 14584
rect 42208 14656 42408 14808
rect 42208 14656 42408 14808
rect 44152 14880 44352 15032
rect 44152 14880 44352 15032
rect 46096 15104 46296 15256
rect 46096 15104 46296 15256
rect 48040 15328 48240 15480
rect 48040 15328 48240 15480
rect 2436 2640 2608 2716
rect 2608 2640 4380 2716
rect 2608 2640 6324 2716
rect 2608 2640 8268 2716
rect 2608 2640 10212 2716
rect 2608 2640 12156 2716
rect 2608 2640 14100 2716
rect 2608 2640 16044 2716
rect 2608 2640 17988 2716
rect 2608 2640 19932 2716
rect 2608 2640 21876 2716
rect 2608 2640 23820 2716
rect 2608 2640 25764 2716
rect 2608 2640 27708 2716
rect 2608 2640 29652 2716
rect 2608 2640 31596 2716
rect 2608 2640 33540 2716
rect 2608 2640 35484 2716
rect 2608 2640 37428 2716
rect 2608 2640 39372 2716
rect 2608 2640 41316 2716
rect 2608 2640 43260 2716
rect 2608 2640 45204 2716
rect 2608 2640 47148 2716
rect 2608 2640 49092 2716
rect 2608 2640 2684 2716
rect 0 2640 216 2728
rect 0 2640 216 2728
rect 2188 2640 2436 2716
rect 108 2640 2188 2716
rect 2188 2640 2264 2716
rect 0 12740 48600 12892
rect 784 12740 25224 12816
rect 784 12740 24300 12816
rect 784 12740 860 12816
rect 0 924 48600 1076
rect 784 924 25224 1000
rect 784 924 24300 1000
rect 784 924 860 1000
<< m3 >>
rect 2398 924 2474 5896
rect 4342 924 4418 5896
rect 6286 924 6362 5896
rect 8230 924 8306 5896
rect 10174 924 10250 5896
rect 12118 924 12194 5896
rect 14062 924 14138 5896
rect 16006 924 16082 5896
rect 17950 924 18026 5896
rect 19894 924 19970 5896
rect 21838 924 21914 5896
rect 23782 924 23858 5896
rect 25726 924 25802 5896
rect 27670 924 27746 5896
rect 29614 924 29690 5896
rect 31558 924 31634 5896
rect 33502 924 33578 5896
rect 35446 924 35522 5896
rect 36446 924 36522 8888
rect 37390 924 37466 5896
rect 39334 924 39410 5896
rect 41278 924 41354 5896
rect 43222 924 43298 5896
rect 45166 924 45242 5896
rect 47110 924 47186 5896
rect 49054 924 49130 5896
<< m1 >>
rect 2406 8976 2466 12892
rect 4350 8976 4410 12892
rect 6294 8976 6354 12892
rect 8238 8976 8298 12892
rect 10182 8976 10242 12892
rect 12126 8976 12186 12892
rect 14070 8976 14130 12892
rect 16014 8976 16074 12892
rect 17958 8976 18018 12892
rect 19902 8976 19962 12892
rect 21846 8976 21906 12892
rect 23790 8976 23850 12892
rect 25734 8976 25794 12892
rect 27678 8976 27738 12892
rect 29622 8976 29682 12892
rect 31566 8976 31626 12892
rect 33510 8976 33570 12892
rect 35454 8976 35514 12892
rect 37398 8976 37458 12892
rect 39342 8976 39402 12892
rect 41286 8976 41346 12892
rect 43230 8976 43290 12892
rect 45174 8976 45234 12892
rect 47118 8976 47178 12892
rect 49062 8976 49122 12892
rect 1396 8800 1572 13920
rect 3340 8800 3516 13920
rect 5284 8800 5460 13920
rect 7228 8800 7404 13920
rect 11116 8800 11292 13920
rect 13060 8800 13236 13920
rect 15004 8800 15180 13920
rect 16948 8800 17124 13920
rect 18892 8800 19068 13920
rect 20836 8800 21012 13920
rect 22780 8800 22956 13920
rect 24724 8800 24900 13920
rect 28612 8800 28788 13920
rect 30556 8800 30732 13920
rect 32500 8800 32676 13920
rect 34444 8800 34620 13920
rect 9172 8800 9348 14360
rect 26668 8800 26844 14360
rect 40276 8800 40452 14584
rect 42220 8800 42396 14808
rect 44164 8800 44340 15032
rect 46108 8800 46284 15256
rect 48052 8800 48228 15480
<< locali >>
rect 49812 336 50112 13480
rect 336 336 50112 636
rect 336 13180 50112 13480
rect 336 336 636 13480
rect 49812 336 50112 13480
rect 816 336 1032 1584
rect 816 336 1032 2376
rect 816 336 1032 5544
rect 816 336 1032 8712
rect 816 336 1032 11880
rect 2760 336 2976 1584
rect 2760 336 2976 2376
rect 2760 336 2976 5544
rect 2760 336 2976 8712
rect 2760 336 2976 11880
rect 4704 336 4920 1584
rect 4704 336 4920 2376
rect 4704 336 4920 5544
rect 4704 336 4920 8712
rect 4704 336 4920 11880
rect 6648 336 6864 1584
rect 6648 336 6864 2376
rect 6648 336 6864 5544
rect 6648 336 6864 8712
rect 6648 336 6864 11880
rect 8592 336 8808 1584
rect 8592 336 8808 2376
rect 8592 336 8808 5544
rect 8592 336 8808 8712
rect 8592 336 8808 11880
rect 10536 336 10752 1584
rect 10536 336 10752 2376
rect 10536 336 10752 5544
rect 10536 336 10752 8712
rect 10536 336 10752 11880
rect 12480 336 12696 1584
rect 12480 336 12696 2376
rect 12480 336 12696 5544
rect 12480 336 12696 8712
rect 12480 336 12696 11880
rect 14424 336 14640 1584
rect 14424 336 14640 2376
rect 14424 336 14640 5544
rect 14424 336 14640 8712
rect 14424 336 14640 11880
rect 16368 336 16584 1584
rect 16368 336 16584 2376
rect 16368 336 16584 5544
rect 16368 336 16584 8712
rect 16368 336 16584 11880
rect 18312 336 18528 1584
rect 18312 336 18528 2376
rect 18312 336 18528 5544
rect 18312 336 18528 8712
rect 18312 336 18528 11880
rect 20256 336 20472 1584
rect 20256 336 20472 2376
rect 20256 336 20472 5544
rect 20256 336 20472 8712
rect 20256 336 20472 11880
rect 22200 336 22416 1584
rect 22200 336 22416 2376
rect 22200 336 22416 5544
rect 22200 336 22416 8712
rect 22200 336 22416 11880
rect 24144 336 24360 1584
rect 24144 336 24360 2376
rect 24144 336 24360 5544
rect 24144 336 24360 8712
rect 24144 336 24360 11880
rect 26088 336 26304 1584
rect 26088 336 26304 2376
rect 26088 336 26304 5544
rect 26088 336 26304 8712
rect 26088 336 26304 11880
rect 28032 336 28248 1584
rect 28032 336 28248 2376
rect 28032 336 28248 5544
rect 28032 336 28248 8712
rect 28032 336 28248 11880
rect 29976 336 30192 1584
rect 29976 336 30192 2376
rect 29976 336 30192 5544
rect 29976 336 30192 8712
rect 29976 336 30192 11880
rect 31920 336 32136 1584
rect 31920 336 32136 2376
rect 31920 336 32136 5544
rect 31920 336 32136 8712
rect 31920 336 32136 11880
rect 33864 336 34080 1584
rect 33864 336 34080 2376
rect 33864 336 34080 5544
rect 33864 336 34080 8712
rect 33864 336 34080 11880
rect 35808 336 36024 1584
rect 35808 336 36024 2376
rect 35808 336 36024 5544
rect 35808 336 36024 8712
rect 35808 336 36024 11880
rect 37752 336 37968 1584
rect 37752 336 37968 2376
rect 37752 336 37968 5544
rect 37752 336 37968 8712
rect 37752 336 37968 11880
rect 39696 336 39912 1584
rect 39696 336 39912 2376
rect 39696 336 39912 5544
rect 39696 336 39912 8712
rect 39696 336 39912 11880
rect 41640 336 41856 1584
rect 41640 336 41856 2376
rect 41640 336 41856 5544
rect 41640 336 41856 8712
rect 41640 336 41856 11880
rect 43584 336 43800 1584
rect 43584 336 43800 2376
rect 43584 336 43800 5544
rect 43584 336 43800 8712
rect 43584 336 43800 11880
rect 45528 336 45744 1584
rect 45528 336 45744 2376
rect 45528 336 45744 5544
rect 45528 336 45744 8712
rect 45528 336 45744 11880
rect 47472 336 47688 1584
rect 47472 336 47688 2376
rect 47472 336 47688 5544
rect 47472 336 47688 8712
rect 47472 336 47688 11880
rect 16 16 50432 128
rect 128 16 50320 128
rect 128 15688 50320 15800
rect 16 15688 50432 15800
rect 16 128 128 15688
rect 16 16 128 15800
rect 50320 128 50432 15688
rect 50320 16 50432 15800
rect 16 16 50432 128
rect 38328 8800 39048 8888
<< ptapc >>
rect 144 32 224 112
rect 224 32 304 112
rect 304 32 384 112
rect 384 32 464 112
rect 464 32 544 112
rect 544 32 624 112
rect 624 32 704 112
rect 704 32 784 112
rect 784 32 864 112
rect 864 32 944 112
rect 944 32 1024 112
rect 1024 32 1104 112
rect 1104 32 1184 112
rect 1184 32 1264 112
rect 1264 32 1344 112
rect 1344 32 1424 112
rect 1424 32 1504 112
rect 1504 32 1584 112
rect 1584 32 1664 112
rect 1664 32 1744 112
rect 1744 32 1824 112
rect 1824 32 1904 112
rect 1904 32 1984 112
rect 1984 32 2064 112
rect 2064 32 2144 112
rect 2144 32 2224 112
rect 2224 32 2304 112
rect 2304 32 2384 112
rect 2384 32 2464 112
rect 2464 32 2544 112
rect 2544 32 2624 112
rect 2624 32 2704 112
rect 2704 32 2784 112
rect 2784 32 2864 112
rect 2864 32 2944 112
rect 2944 32 3024 112
rect 3024 32 3104 112
rect 3104 32 3184 112
rect 3184 32 3264 112
rect 3264 32 3344 112
rect 3344 32 3424 112
rect 3424 32 3504 112
rect 3504 32 3584 112
rect 3584 32 3664 112
rect 3664 32 3744 112
rect 3744 32 3824 112
rect 3824 32 3904 112
rect 3904 32 3984 112
rect 3984 32 4064 112
rect 4064 32 4144 112
rect 4144 32 4224 112
rect 4224 32 4304 112
rect 4304 32 4384 112
rect 4384 32 4464 112
rect 4464 32 4544 112
rect 4544 32 4624 112
rect 4624 32 4704 112
rect 4704 32 4784 112
rect 4784 32 4864 112
rect 4864 32 4944 112
rect 4944 32 5024 112
rect 5024 32 5104 112
rect 5104 32 5184 112
rect 5184 32 5264 112
rect 5264 32 5344 112
rect 5344 32 5424 112
rect 5424 32 5504 112
rect 5504 32 5584 112
rect 5584 32 5664 112
rect 5664 32 5744 112
rect 5744 32 5824 112
rect 5824 32 5904 112
rect 5904 32 5984 112
rect 5984 32 6064 112
rect 6064 32 6144 112
rect 6144 32 6224 112
rect 6224 32 6304 112
rect 6304 32 6384 112
rect 6384 32 6464 112
rect 6464 32 6544 112
rect 6544 32 6624 112
rect 6624 32 6704 112
rect 6704 32 6784 112
rect 6784 32 6864 112
rect 6864 32 6944 112
rect 6944 32 7024 112
rect 7024 32 7104 112
rect 7104 32 7184 112
rect 7184 32 7264 112
rect 7264 32 7344 112
rect 7344 32 7424 112
rect 7424 32 7504 112
rect 7504 32 7584 112
rect 7584 32 7664 112
rect 7664 32 7744 112
rect 7744 32 7824 112
rect 7824 32 7904 112
rect 7904 32 7984 112
rect 7984 32 8064 112
rect 8064 32 8144 112
rect 8144 32 8224 112
rect 8224 32 8304 112
rect 8304 32 8384 112
rect 8384 32 8464 112
rect 8464 32 8544 112
rect 8544 32 8624 112
rect 8624 32 8704 112
rect 8704 32 8784 112
rect 8784 32 8864 112
rect 8864 32 8944 112
rect 8944 32 9024 112
rect 9024 32 9104 112
rect 9104 32 9184 112
rect 9184 32 9264 112
rect 9264 32 9344 112
rect 9344 32 9424 112
rect 9424 32 9504 112
rect 9504 32 9584 112
rect 9584 32 9664 112
rect 9664 32 9744 112
rect 9744 32 9824 112
rect 9824 32 9904 112
rect 9904 32 9984 112
rect 9984 32 10064 112
rect 10064 32 10144 112
rect 10144 32 10224 112
rect 10224 32 10304 112
rect 10304 32 10384 112
rect 10384 32 10464 112
rect 10464 32 10544 112
rect 10544 32 10624 112
rect 10624 32 10704 112
rect 10704 32 10784 112
rect 10784 32 10864 112
rect 10864 32 10944 112
rect 10944 32 11024 112
rect 11024 32 11104 112
rect 11104 32 11184 112
rect 11184 32 11264 112
rect 11264 32 11344 112
rect 11344 32 11424 112
rect 11424 32 11504 112
rect 11504 32 11584 112
rect 11584 32 11664 112
rect 11664 32 11744 112
rect 11744 32 11824 112
rect 11824 32 11904 112
rect 11904 32 11984 112
rect 11984 32 12064 112
rect 12064 32 12144 112
rect 12144 32 12224 112
rect 12224 32 12304 112
rect 12304 32 12384 112
rect 12384 32 12464 112
rect 12464 32 12544 112
rect 12544 32 12624 112
rect 12624 32 12704 112
rect 12704 32 12784 112
rect 12784 32 12864 112
rect 12864 32 12944 112
rect 12944 32 13024 112
rect 13024 32 13104 112
rect 13104 32 13184 112
rect 13184 32 13264 112
rect 13264 32 13344 112
rect 13344 32 13424 112
rect 13424 32 13504 112
rect 13504 32 13584 112
rect 13584 32 13664 112
rect 13664 32 13744 112
rect 13744 32 13824 112
rect 13824 32 13904 112
rect 13904 32 13984 112
rect 13984 32 14064 112
rect 14064 32 14144 112
rect 14144 32 14224 112
rect 14224 32 14304 112
rect 14304 32 14384 112
rect 14384 32 14464 112
rect 14464 32 14544 112
rect 14544 32 14624 112
rect 14624 32 14704 112
rect 14704 32 14784 112
rect 14784 32 14864 112
rect 14864 32 14944 112
rect 14944 32 15024 112
rect 15024 32 15104 112
rect 15104 32 15184 112
rect 15184 32 15264 112
rect 15264 32 15344 112
rect 15344 32 15424 112
rect 15424 32 15504 112
rect 15504 32 15584 112
rect 15584 32 15664 112
rect 15664 32 15744 112
rect 15744 32 15824 112
rect 15824 32 15904 112
rect 15904 32 15984 112
rect 15984 32 16064 112
rect 16064 32 16144 112
rect 16144 32 16224 112
rect 16224 32 16304 112
rect 16304 32 16384 112
rect 16384 32 16464 112
rect 16464 32 16544 112
rect 16544 32 16624 112
rect 16624 32 16704 112
rect 16704 32 16784 112
rect 16784 32 16864 112
rect 16864 32 16944 112
rect 16944 32 17024 112
rect 17024 32 17104 112
rect 17104 32 17184 112
rect 17184 32 17264 112
rect 17264 32 17344 112
rect 17344 32 17424 112
rect 17424 32 17504 112
rect 17504 32 17584 112
rect 17584 32 17664 112
rect 17664 32 17744 112
rect 17744 32 17824 112
rect 17824 32 17904 112
rect 17904 32 17984 112
rect 17984 32 18064 112
rect 18064 32 18144 112
rect 18144 32 18224 112
rect 18224 32 18304 112
rect 18304 32 18384 112
rect 18384 32 18464 112
rect 18464 32 18544 112
rect 18544 32 18624 112
rect 18624 32 18704 112
rect 18704 32 18784 112
rect 18784 32 18864 112
rect 18864 32 18944 112
rect 18944 32 19024 112
rect 19024 32 19104 112
rect 19104 32 19184 112
rect 19184 32 19264 112
rect 19264 32 19344 112
rect 19344 32 19424 112
rect 19424 32 19504 112
rect 19504 32 19584 112
rect 19584 32 19664 112
rect 19664 32 19744 112
rect 19744 32 19824 112
rect 19824 32 19904 112
rect 19904 32 19984 112
rect 19984 32 20064 112
rect 20064 32 20144 112
rect 20144 32 20224 112
rect 20224 32 20304 112
rect 20304 32 20384 112
rect 20384 32 20464 112
rect 20464 32 20544 112
rect 20544 32 20624 112
rect 20624 32 20704 112
rect 20704 32 20784 112
rect 20784 32 20864 112
rect 20864 32 20944 112
rect 20944 32 21024 112
rect 21024 32 21104 112
rect 21104 32 21184 112
rect 21184 32 21264 112
rect 21264 32 21344 112
rect 21344 32 21424 112
rect 21424 32 21504 112
rect 21504 32 21584 112
rect 21584 32 21664 112
rect 21664 32 21744 112
rect 21744 32 21824 112
rect 21824 32 21904 112
rect 21904 32 21984 112
rect 21984 32 22064 112
rect 22064 32 22144 112
rect 22144 32 22224 112
rect 22224 32 22304 112
rect 22304 32 22384 112
rect 22384 32 22464 112
rect 22464 32 22544 112
rect 22544 32 22624 112
rect 22624 32 22704 112
rect 22704 32 22784 112
rect 22784 32 22864 112
rect 22864 32 22944 112
rect 22944 32 23024 112
rect 23024 32 23104 112
rect 23104 32 23184 112
rect 23184 32 23264 112
rect 23264 32 23344 112
rect 23344 32 23424 112
rect 23424 32 23504 112
rect 23504 32 23584 112
rect 23584 32 23664 112
rect 23664 32 23744 112
rect 23744 32 23824 112
rect 23824 32 23904 112
rect 23904 32 23984 112
rect 23984 32 24064 112
rect 24064 32 24144 112
rect 24144 32 24224 112
rect 24224 32 24304 112
rect 24304 32 24384 112
rect 24384 32 24464 112
rect 24464 32 24544 112
rect 24544 32 24624 112
rect 24624 32 24704 112
rect 24704 32 24784 112
rect 24784 32 24864 112
rect 24864 32 24944 112
rect 24944 32 25024 112
rect 25024 32 25104 112
rect 25104 32 25184 112
rect 25184 32 25264 112
rect 25264 32 25344 112
rect 25344 32 25424 112
rect 25424 32 25504 112
rect 25504 32 25584 112
rect 25584 32 25664 112
rect 25664 32 25744 112
rect 25744 32 25824 112
rect 25824 32 25904 112
rect 25904 32 25984 112
rect 25984 32 26064 112
rect 26064 32 26144 112
rect 26144 32 26224 112
rect 26224 32 26304 112
rect 26304 32 26384 112
rect 26384 32 26464 112
rect 26464 32 26544 112
rect 26544 32 26624 112
rect 26624 32 26704 112
rect 26704 32 26784 112
rect 26784 32 26864 112
rect 26864 32 26944 112
rect 26944 32 27024 112
rect 27024 32 27104 112
rect 27104 32 27184 112
rect 27184 32 27264 112
rect 27264 32 27344 112
rect 27344 32 27424 112
rect 27424 32 27504 112
rect 27504 32 27584 112
rect 27584 32 27664 112
rect 27664 32 27744 112
rect 27744 32 27824 112
rect 27824 32 27904 112
rect 27904 32 27984 112
rect 27984 32 28064 112
rect 28064 32 28144 112
rect 28144 32 28224 112
rect 28224 32 28304 112
rect 28304 32 28384 112
rect 28384 32 28464 112
rect 28464 32 28544 112
rect 28544 32 28624 112
rect 28624 32 28704 112
rect 28704 32 28784 112
rect 28784 32 28864 112
rect 28864 32 28944 112
rect 28944 32 29024 112
rect 29024 32 29104 112
rect 29104 32 29184 112
rect 29184 32 29264 112
rect 29264 32 29344 112
rect 29344 32 29424 112
rect 29424 32 29504 112
rect 29504 32 29584 112
rect 29584 32 29664 112
rect 29664 32 29744 112
rect 29744 32 29824 112
rect 29824 32 29904 112
rect 29904 32 29984 112
rect 29984 32 30064 112
rect 30064 32 30144 112
rect 30144 32 30224 112
rect 30224 32 30304 112
rect 30304 32 30384 112
rect 30384 32 30464 112
rect 30464 32 30544 112
rect 30544 32 30624 112
rect 30624 32 30704 112
rect 30704 32 30784 112
rect 30784 32 30864 112
rect 30864 32 30944 112
rect 30944 32 31024 112
rect 31024 32 31104 112
rect 31104 32 31184 112
rect 31184 32 31264 112
rect 31264 32 31344 112
rect 31344 32 31424 112
rect 31424 32 31504 112
rect 31504 32 31584 112
rect 31584 32 31664 112
rect 31664 32 31744 112
rect 31744 32 31824 112
rect 31824 32 31904 112
rect 31904 32 31984 112
rect 31984 32 32064 112
rect 32064 32 32144 112
rect 32144 32 32224 112
rect 32224 32 32304 112
rect 32304 32 32384 112
rect 32384 32 32464 112
rect 32464 32 32544 112
rect 32544 32 32624 112
rect 32624 32 32704 112
rect 32704 32 32784 112
rect 32784 32 32864 112
rect 32864 32 32944 112
rect 32944 32 33024 112
rect 33024 32 33104 112
rect 33104 32 33184 112
rect 33184 32 33264 112
rect 33264 32 33344 112
rect 33344 32 33424 112
rect 33424 32 33504 112
rect 33504 32 33584 112
rect 33584 32 33664 112
rect 33664 32 33744 112
rect 33744 32 33824 112
rect 33824 32 33904 112
rect 33904 32 33984 112
rect 33984 32 34064 112
rect 34064 32 34144 112
rect 34144 32 34224 112
rect 34224 32 34304 112
rect 34304 32 34384 112
rect 34384 32 34464 112
rect 34464 32 34544 112
rect 34544 32 34624 112
rect 34624 32 34704 112
rect 34704 32 34784 112
rect 34784 32 34864 112
rect 34864 32 34944 112
rect 34944 32 35024 112
rect 35024 32 35104 112
rect 35104 32 35184 112
rect 35184 32 35264 112
rect 35264 32 35344 112
rect 35344 32 35424 112
rect 35424 32 35504 112
rect 35504 32 35584 112
rect 35584 32 35664 112
rect 35664 32 35744 112
rect 35744 32 35824 112
rect 35824 32 35904 112
rect 35904 32 35984 112
rect 35984 32 36064 112
rect 36064 32 36144 112
rect 36144 32 36224 112
rect 36224 32 36304 112
rect 36304 32 36384 112
rect 36384 32 36464 112
rect 36464 32 36544 112
rect 36544 32 36624 112
rect 36624 32 36704 112
rect 36704 32 36784 112
rect 36784 32 36864 112
rect 36864 32 36944 112
rect 36944 32 37024 112
rect 37024 32 37104 112
rect 37104 32 37184 112
rect 37184 32 37264 112
rect 37264 32 37344 112
rect 37344 32 37424 112
rect 37424 32 37504 112
rect 37504 32 37584 112
rect 37584 32 37664 112
rect 37664 32 37744 112
rect 37744 32 37824 112
rect 37824 32 37904 112
rect 37904 32 37984 112
rect 37984 32 38064 112
rect 38064 32 38144 112
rect 38144 32 38224 112
rect 38224 32 38304 112
rect 38304 32 38384 112
rect 38384 32 38464 112
rect 38464 32 38544 112
rect 38544 32 38624 112
rect 38624 32 38704 112
rect 38704 32 38784 112
rect 38784 32 38864 112
rect 38864 32 38944 112
rect 38944 32 39024 112
rect 39024 32 39104 112
rect 39104 32 39184 112
rect 39184 32 39264 112
rect 39264 32 39344 112
rect 39344 32 39424 112
rect 39424 32 39504 112
rect 39504 32 39584 112
rect 39584 32 39664 112
rect 39664 32 39744 112
rect 39744 32 39824 112
rect 39824 32 39904 112
rect 39904 32 39984 112
rect 39984 32 40064 112
rect 40064 32 40144 112
rect 40144 32 40224 112
rect 40224 32 40304 112
rect 40304 32 40384 112
rect 40384 32 40464 112
rect 40464 32 40544 112
rect 40544 32 40624 112
rect 40624 32 40704 112
rect 40704 32 40784 112
rect 40784 32 40864 112
rect 40864 32 40944 112
rect 40944 32 41024 112
rect 41024 32 41104 112
rect 41104 32 41184 112
rect 41184 32 41264 112
rect 41264 32 41344 112
rect 41344 32 41424 112
rect 41424 32 41504 112
rect 41504 32 41584 112
rect 41584 32 41664 112
rect 41664 32 41744 112
rect 41744 32 41824 112
rect 41824 32 41904 112
rect 41904 32 41984 112
rect 41984 32 42064 112
rect 42064 32 42144 112
rect 42144 32 42224 112
rect 42224 32 42304 112
rect 42304 32 42384 112
rect 42384 32 42464 112
rect 42464 32 42544 112
rect 42544 32 42624 112
rect 42624 32 42704 112
rect 42704 32 42784 112
rect 42784 32 42864 112
rect 42864 32 42944 112
rect 42944 32 43024 112
rect 43024 32 43104 112
rect 43104 32 43184 112
rect 43184 32 43264 112
rect 43264 32 43344 112
rect 43344 32 43424 112
rect 43424 32 43504 112
rect 43504 32 43584 112
rect 43584 32 43664 112
rect 43664 32 43744 112
rect 43744 32 43824 112
rect 43824 32 43904 112
rect 43904 32 43984 112
rect 43984 32 44064 112
rect 44064 32 44144 112
rect 44144 32 44224 112
rect 44224 32 44304 112
rect 44304 32 44384 112
rect 44384 32 44464 112
rect 44464 32 44544 112
rect 44544 32 44624 112
rect 44624 32 44704 112
rect 44704 32 44784 112
rect 44784 32 44864 112
rect 44864 32 44944 112
rect 44944 32 45024 112
rect 45024 32 45104 112
rect 45104 32 45184 112
rect 45184 32 45264 112
rect 45264 32 45344 112
rect 45344 32 45424 112
rect 45424 32 45504 112
rect 45504 32 45584 112
rect 45584 32 45664 112
rect 45664 32 45744 112
rect 45744 32 45824 112
rect 45824 32 45904 112
rect 45904 32 45984 112
rect 45984 32 46064 112
rect 46064 32 46144 112
rect 46144 32 46224 112
rect 46224 32 46304 112
rect 46304 32 46384 112
rect 46384 32 46464 112
rect 46464 32 46544 112
rect 46544 32 46624 112
rect 46624 32 46704 112
rect 46704 32 46784 112
rect 46784 32 46864 112
rect 46864 32 46944 112
rect 46944 32 47024 112
rect 47024 32 47104 112
rect 47104 32 47184 112
rect 47184 32 47264 112
rect 47264 32 47344 112
rect 47344 32 47424 112
rect 47424 32 47504 112
rect 47504 32 47584 112
rect 47584 32 47664 112
rect 47664 32 47744 112
rect 47744 32 47824 112
rect 47824 32 47904 112
rect 47904 32 47984 112
rect 47984 32 48064 112
rect 48064 32 48144 112
rect 48144 32 48224 112
rect 48224 32 48304 112
rect 48304 32 48384 112
rect 48384 32 48464 112
rect 48464 32 48544 112
rect 48544 32 48624 112
rect 48624 32 48704 112
rect 48704 32 48784 112
rect 48784 32 48864 112
rect 48864 32 48944 112
rect 48944 32 49024 112
rect 49024 32 49104 112
rect 49104 32 49184 112
rect 49184 32 49264 112
rect 49264 32 49344 112
rect 49344 32 49424 112
rect 49424 32 49504 112
rect 49504 32 49584 112
rect 49584 32 49664 112
rect 49664 32 49744 112
rect 49744 32 49824 112
rect 49824 32 49904 112
rect 49904 32 49984 112
rect 49984 32 50064 112
rect 50064 32 50144 112
rect 50144 32 50224 112
rect 50224 32 50304 112
rect 144 15704 224 15784
rect 224 15704 304 15784
rect 304 15704 384 15784
rect 384 15704 464 15784
rect 464 15704 544 15784
rect 544 15704 624 15784
rect 624 15704 704 15784
rect 704 15704 784 15784
rect 784 15704 864 15784
rect 864 15704 944 15784
rect 944 15704 1024 15784
rect 1024 15704 1104 15784
rect 1104 15704 1184 15784
rect 1184 15704 1264 15784
rect 1264 15704 1344 15784
rect 1344 15704 1424 15784
rect 1424 15704 1504 15784
rect 1504 15704 1584 15784
rect 1584 15704 1664 15784
rect 1664 15704 1744 15784
rect 1744 15704 1824 15784
rect 1824 15704 1904 15784
rect 1904 15704 1984 15784
rect 1984 15704 2064 15784
rect 2064 15704 2144 15784
rect 2144 15704 2224 15784
rect 2224 15704 2304 15784
rect 2304 15704 2384 15784
rect 2384 15704 2464 15784
rect 2464 15704 2544 15784
rect 2544 15704 2624 15784
rect 2624 15704 2704 15784
rect 2704 15704 2784 15784
rect 2784 15704 2864 15784
rect 2864 15704 2944 15784
rect 2944 15704 3024 15784
rect 3024 15704 3104 15784
rect 3104 15704 3184 15784
rect 3184 15704 3264 15784
rect 3264 15704 3344 15784
rect 3344 15704 3424 15784
rect 3424 15704 3504 15784
rect 3504 15704 3584 15784
rect 3584 15704 3664 15784
rect 3664 15704 3744 15784
rect 3744 15704 3824 15784
rect 3824 15704 3904 15784
rect 3904 15704 3984 15784
rect 3984 15704 4064 15784
rect 4064 15704 4144 15784
rect 4144 15704 4224 15784
rect 4224 15704 4304 15784
rect 4304 15704 4384 15784
rect 4384 15704 4464 15784
rect 4464 15704 4544 15784
rect 4544 15704 4624 15784
rect 4624 15704 4704 15784
rect 4704 15704 4784 15784
rect 4784 15704 4864 15784
rect 4864 15704 4944 15784
rect 4944 15704 5024 15784
rect 5024 15704 5104 15784
rect 5104 15704 5184 15784
rect 5184 15704 5264 15784
rect 5264 15704 5344 15784
rect 5344 15704 5424 15784
rect 5424 15704 5504 15784
rect 5504 15704 5584 15784
rect 5584 15704 5664 15784
rect 5664 15704 5744 15784
rect 5744 15704 5824 15784
rect 5824 15704 5904 15784
rect 5904 15704 5984 15784
rect 5984 15704 6064 15784
rect 6064 15704 6144 15784
rect 6144 15704 6224 15784
rect 6224 15704 6304 15784
rect 6304 15704 6384 15784
rect 6384 15704 6464 15784
rect 6464 15704 6544 15784
rect 6544 15704 6624 15784
rect 6624 15704 6704 15784
rect 6704 15704 6784 15784
rect 6784 15704 6864 15784
rect 6864 15704 6944 15784
rect 6944 15704 7024 15784
rect 7024 15704 7104 15784
rect 7104 15704 7184 15784
rect 7184 15704 7264 15784
rect 7264 15704 7344 15784
rect 7344 15704 7424 15784
rect 7424 15704 7504 15784
rect 7504 15704 7584 15784
rect 7584 15704 7664 15784
rect 7664 15704 7744 15784
rect 7744 15704 7824 15784
rect 7824 15704 7904 15784
rect 7904 15704 7984 15784
rect 7984 15704 8064 15784
rect 8064 15704 8144 15784
rect 8144 15704 8224 15784
rect 8224 15704 8304 15784
rect 8304 15704 8384 15784
rect 8384 15704 8464 15784
rect 8464 15704 8544 15784
rect 8544 15704 8624 15784
rect 8624 15704 8704 15784
rect 8704 15704 8784 15784
rect 8784 15704 8864 15784
rect 8864 15704 8944 15784
rect 8944 15704 9024 15784
rect 9024 15704 9104 15784
rect 9104 15704 9184 15784
rect 9184 15704 9264 15784
rect 9264 15704 9344 15784
rect 9344 15704 9424 15784
rect 9424 15704 9504 15784
rect 9504 15704 9584 15784
rect 9584 15704 9664 15784
rect 9664 15704 9744 15784
rect 9744 15704 9824 15784
rect 9824 15704 9904 15784
rect 9904 15704 9984 15784
rect 9984 15704 10064 15784
rect 10064 15704 10144 15784
rect 10144 15704 10224 15784
rect 10224 15704 10304 15784
rect 10304 15704 10384 15784
rect 10384 15704 10464 15784
rect 10464 15704 10544 15784
rect 10544 15704 10624 15784
rect 10624 15704 10704 15784
rect 10704 15704 10784 15784
rect 10784 15704 10864 15784
rect 10864 15704 10944 15784
rect 10944 15704 11024 15784
rect 11024 15704 11104 15784
rect 11104 15704 11184 15784
rect 11184 15704 11264 15784
rect 11264 15704 11344 15784
rect 11344 15704 11424 15784
rect 11424 15704 11504 15784
rect 11504 15704 11584 15784
rect 11584 15704 11664 15784
rect 11664 15704 11744 15784
rect 11744 15704 11824 15784
rect 11824 15704 11904 15784
rect 11904 15704 11984 15784
rect 11984 15704 12064 15784
rect 12064 15704 12144 15784
rect 12144 15704 12224 15784
rect 12224 15704 12304 15784
rect 12304 15704 12384 15784
rect 12384 15704 12464 15784
rect 12464 15704 12544 15784
rect 12544 15704 12624 15784
rect 12624 15704 12704 15784
rect 12704 15704 12784 15784
rect 12784 15704 12864 15784
rect 12864 15704 12944 15784
rect 12944 15704 13024 15784
rect 13024 15704 13104 15784
rect 13104 15704 13184 15784
rect 13184 15704 13264 15784
rect 13264 15704 13344 15784
rect 13344 15704 13424 15784
rect 13424 15704 13504 15784
rect 13504 15704 13584 15784
rect 13584 15704 13664 15784
rect 13664 15704 13744 15784
rect 13744 15704 13824 15784
rect 13824 15704 13904 15784
rect 13904 15704 13984 15784
rect 13984 15704 14064 15784
rect 14064 15704 14144 15784
rect 14144 15704 14224 15784
rect 14224 15704 14304 15784
rect 14304 15704 14384 15784
rect 14384 15704 14464 15784
rect 14464 15704 14544 15784
rect 14544 15704 14624 15784
rect 14624 15704 14704 15784
rect 14704 15704 14784 15784
rect 14784 15704 14864 15784
rect 14864 15704 14944 15784
rect 14944 15704 15024 15784
rect 15024 15704 15104 15784
rect 15104 15704 15184 15784
rect 15184 15704 15264 15784
rect 15264 15704 15344 15784
rect 15344 15704 15424 15784
rect 15424 15704 15504 15784
rect 15504 15704 15584 15784
rect 15584 15704 15664 15784
rect 15664 15704 15744 15784
rect 15744 15704 15824 15784
rect 15824 15704 15904 15784
rect 15904 15704 15984 15784
rect 15984 15704 16064 15784
rect 16064 15704 16144 15784
rect 16144 15704 16224 15784
rect 16224 15704 16304 15784
rect 16304 15704 16384 15784
rect 16384 15704 16464 15784
rect 16464 15704 16544 15784
rect 16544 15704 16624 15784
rect 16624 15704 16704 15784
rect 16704 15704 16784 15784
rect 16784 15704 16864 15784
rect 16864 15704 16944 15784
rect 16944 15704 17024 15784
rect 17024 15704 17104 15784
rect 17104 15704 17184 15784
rect 17184 15704 17264 15784
rect 17264 15704 17344 15784
rect 17344 15704 17424 15784
rect 17424 15704 17504 15784
rect 17504 15704 17584 15784
rect 17584 15704 17664 15784
rect 17664 15704 17744 15784
rect 17744 15704 17824 15784
rect 17824 15704 17904 15784
rect 17904 15704 17984 15784
rect 17984 15704 18064 15784
rect 18064 15704 18144 15784
rect 18144 15704 18224 15784
rect 18224 15704 18304 15784
rect 18304 15704 18384 15784
rect 18384 15704 18464 15784
rect 18464 15704 18544 15784
rect 18544 15704 18624 15784
rect 18624 15704 18704 15784
rect 18704 15704 18784 15784
rect 18784 15704 18864 15784
rect 18864 15704 18944 15784
rect 18944 15704 19024 15784
rect 19024 15704 19104 15784
rect 19104 15704 19184 15784
rect 19184 15704 19264 15784
rect 19264 15704 19344 15784
rect 19344 15704 19424 15784
rect 19424 15704 19504 15784
rect 19504 15704 19584 15784
rect 19584 15704 19664 15784
rect 19664 15704 19744 15784
rect 19744 15704 19824 15784
rect 19824 15704 19904 15784
rect 19904 15704 19984 15784
rect 19984 15704 20064 15784
rect 20064 15704 20144 15784
rect 20144 15704 20224 15784
rect 20224 15704 20304 15784
rect 20304 15704 20384 15784
rect 20384 15704 20464 15784
rect 20464 15704 20544 15784
rect 20544 15704 20624 15784
rect 20624 15704 20704 15784
rect 20704 15704 20784 15784
rect 20784 15704 20864 15784
rect 20864 15704 20944 15784
rect 20944 15704 21024 15784
rect 21024 15704 21104 15784
rect 21104 15704 21184 15784
rect 21184 15704 21264 15784
rect 21264 15704 21344 15784
rect 21344 15704 21424 15784
rect 21424 15704 21504 15784
rect 21504 15704 21584 15784
rect 21584 15704 21664 15784
rect 21664 15704 21744 15784
rect 21744 15704 21824 15784
rect 21824 15704 21904 15784
rect 21904 15704 21984 15784
rect 21984 15704 22064 15784
rect 22064 15704 22144 15784
rect 22144 15704 22224 15784
rect 22224 15704 22304 15784
rect 22304 15704 22384 15784
rect 22384 15704 22464 15784
rect 22464 15704 22544 15784
rect 22544 15704 22624 15784
rect 22624 15704 22704 15784
rect 22704 15704 22784 15784
rect 22784 15704 22864 15784
rect 22864 15704 22944 15784
rect 22944 15704 23024 15784
rect 23024 15704 23104 15784
rect 23104 15704 23184 15784
rect 23184 15704 23264 15784
rect 23264 15704 23344 15784
rect 23344 15704 23424 15784
rect 23424 15704 23504 15784
rect 23504 15704 23584 15784
rect 23584 15704 23664 15784
rect 23664 15704 23744 15784
rect 23744 15704 23824 15784
rect 23824 15704 23904 15784
rect 23904 15704 23984 15784
rect 23984 15704 24064 15784
rect 24064 15704 24144 15784
rect 24144 15704 24224 15784
rect 24224 15704 24304 15784
rect 24304 15704 24384 15784
rect 24384 15704 24464 15784
rect 24464 15704 24544 15784
rect 24544 15704 24624 15784
rect 24624 15704 24704 15784
rect 24704 15704 24784 15784
rect 24784 15704 24864 15784
rect 24864 15704 24944 15784
rect 24944 15704 25024 15784
rect 25024 15704 25104 15784
rect 25104 15704 25184 15784
rect 25184 15704 25264 15784
rect 25264 15704 25344 15784
rect 25344 15704 25424 15784
rect 25424 15704 25504 15784
rect 25504 15704 25584 15784
rect 25584 15704 25664 15784
rect 25664 15704 25744 15784
rect 25744 15704 25824 15784
rect 25824 15704 25904 15784
rect 25904 15704 25984 15784
rect 25984 15704 26064 15784
rect 26064 15704 26144 15784
rect 26144 15704 26224 15784
rect 26224 15704 26304 15784
rect 26304 15704 26384 15784
rect 26384 15704 26464 15784
rect 26464 15704 26544 15784
rect 26544 15704 26624 15784
rect 26624 15704 26704 15784
rect 26704 15704 26784 15784
rect 26784 15704 26864 15784
rect 26864 15704 26944 15784
rect 26944 15704 27024 15784
rect 27024 15704 27104 15784
rect 27104 15704 27184 15784
rect 27184 15704 27264 15784
rect 27264 15704 27344 15784
rect 27344 15704 27424 15784
rect 27424 15704 27504 15784
rect 27504 15704 27584 15784
rect 27584 15704 27664 15784
rect 27664 15704 27744 15784
rect 27744 15704 27824 15784
rect 27824 15704 27904 15784
rect 27904 15704 27984 15784
rect 27984 15704 28064 15784
rect 28064 15704 28144 15784
rect 28144 15704 28224 15784
rect 28224 15704 28304 15784
rect 28304 15704 28384 15784
rect 28384 15704 28464 15784
rect 28464 15704 28544 15784
rect 28544 15704 28624 15784
rect 28624 15704 28704 15784
rect 28704 15704 28784 15784
rect 28784 15704 28864 15784
rect 28864 15704 28944 15784
rect 28944 15704 29024 15784
rect 29024 15704 29104 15784
rect 29104 15704 29184 15784
rect 29184 15704 29264 15784
rect 29264 15704 29344 15784
rect 29344 15704 29424 15784
rect 29424 15704 29504 15784
rect 29504 15704 29584 15784
rect 29584 15704 29664 15784
rect 29664 15704 29744 15784
rect 29744 15704 29824 15784
rect 29824 15704 29904 15784
rect 29904 15704 29984 15784
rect 29984 15704 30064 15784
rect 30064 15704 30144 15784
rect 30144 15704 30224 15784
rect 30224 15704 30304 15784
rect 30304 15704 30384 15784
rect 30384 15704 30464 15784
rect 30464 15704 30544 15784
rect 30544 15704 30624 15784
rect 30624 15704 30704 15784
rect 30704 15704 30784 15784
rect 30784 15704 30864 15784
rect 30864 15704 30944 15784
rect 30944 15704 31024 15784
rect 31024 15704 31104 15784
rect 31104 15704 31184 15784
rect 31184 15704 31264 15784
rect 31264 15704 31344 15784
rect 31344 15704 31424 15784
rect 31424 15704 31504 15784
rect 31504 15704 31584 15784
rect 31584 15704 31664 15784
rect 31664 15704 31744 15784
rect 31744 15704 31824 15784
rect 31824 15704 31904 15784
rect 31904 15704 31984 15784
rect 31984 15704 32064 15784
rect 32064 15704 32144 15784
rect 32144 15704 32224 15784
rect 32224 15704 32304 15784
rect 32304 15704 32384 15784
rect 32384 15704 32464 15784
rect 32464 15704 32544 15784
rect 32544 15704 32624 15784
rect 32624 15704 32704 15784
rect 32704 15704 32784 15784
rect 32784 15704 32864 15784
rect 32864 15704 32944 15784
rect 32944 15704 33024 15784
rect 33024 15704 33104 15784
rect 33104 15704 33184 15784
rect 33184 15704 33264 15784
rect 33264 15704 33344 15784
rect 33344 15704 33424 15784
rect 33424 15704 33504 15784
rect 33504 15704 33584 15784
rect 33584 15704 33664 15784
rect 33664 15704 33744 15784
rect 33744 15704 33824 15784
rect 33824 15704 33904 15784
rect 33904 15704 33984 15784
rect 33984 15704 34064 15784
rect 34064 15704 34144 15784
rect 34144 15704 34224 15784
rect 34224 15704 34304 15784
rect 34304 15704 34384 15784
rect 34384 15704 34464 15784
rect 34464 15704 34544 15784
rect 34544 15704 34624 15784
rect 34624 15704 34704 15784
rect 34704 15704 34784 15784
rect 34784 15704 34864 15784
rect 34864 15704 34944 15784
rect 34944 15704 35024 15784
rect 35024 15704 35104 15784
rect 35104 15704 35184 15784
rect 35184 15704 35264 15784
rect 35264 15704 35344 15784
rect 35344 15704 35424 15784
rect 35424 15704 35504 15784
rect 35504 15704 35584 15784
rect 35584 15704 35664 15784
rect 35664 15704 35744 15784
rect 35744 15704 35824 15784
rect 35824 15704 35904 15784
rect 35904 15704 35984 15784
rect 35984 15704 36064 15784
rect 36064 15704 36144 15784
rect 36144 15704 36224 15784
rect 36224 15704 36304 15784
rect 36304 15704 36384 15784
rect 36384 15704 36464 15784
rect 36464 15704 36544 15784
rect 36544 15704 36624 15784
rect 36624 15704 36704 15784
rect 36704 15704 36784 15784
rect 36784 15704 36864 15784
rect 36864 15704 36944 15784
rect 36944 15704 37024 15784
rect 37024 15704 37104 15784
rect 37104 15704 37184 15784
rect 37184 15704 37264 15784
rect 37264 15704 37344 15784
rect 37344 15704 37424 15784
rect 37424 15704 37504 15784
rect 37504 15704 37584 15784
rect 37584 15704 37664 15784
rect 37664 15704 37744 15784
rect 37744 15704 37824 15784
rect 37824 15704 37904 15784
rect 37904 15704 37984 15784
rect 37984 15704 38064 15784
rect 38064 15704 38144 15784
rect 38144 15704 38224 15784
rect 38224 15704 38304 15784
rect 38304 15704 38384 15784
rect 38384 15704 38464 15784
rect 38464 15704 38544 15784
rect 38544 15704 38624 15784
rect 38624 15704 38704 15784
rect 38704 15704 38784 15784
rect 38784 15704 38864 15784
rect 38864 15704 38944 15784
rect 38944 15704 39024 15784
rect 39024 15704 39104 15784
rect 39104 15704 39184 15784
rect 39184 15704 39264 15784
rect 39264 15704 39344 15784
rect 39344 15704 39424 15784
rect 39424 15704 39504 15784
rect 39504 15704 39584 15784
rect 39584 15704 39664 15784
rect 39664 15704 39744 15784
rect 39744 15704 39824 15784
rect 39824 15704 39904 15784
rect 39904 15704 39984 15784
rect 39984 15704 40064 15784
rect 40064 15704 40144 15784
rect 40144 15704 40224 15784
rect 40224 15704 40304 15784
rect 40304 15704 40384 15784
rect 40384 15704 40464 15784
rect 40464 15704 40544 15784
rect 40544 15704 40624 15784
rect 40624 15704 40704 15784
rect 40704 15704 40784 15784
rect 40784 15704 40864 15784
rect 40864 15704 40944 15784
rect 40944 15704 41024 15784
rect 41024 15704 41104 15784
rect 41104 15704 41184 15784
rect 41184 15704 41264 15784
rect 41264 15704 41344 15784
rect 41344 15704 41424 15784
rect 41424 15704 41504 15784
rect 41504 15704 41584 15784
rect 41584 15704 41664 15784
rect 41664 15704 41744 15784
rect 41744 15704 41824 15784
rect 41824 15704 41904 15784
rect 41904 15704 41984 15784
rect 41984 15704 42064 15784
rect 42064 15704 42144 15784
rect 42144 15704 42224 15784
rect 42224 15704 42304 15784
rect 42304 15704 42384 15784
rect 42384 15704 42464 15784
rect 42464 15704 42544 15784
rect 42544 15704 42624 15784
rect 42624 15704 42704 15784
rect 42704 15704 42784 15784
rect 42784 15704 42864 15784
rect 42864 15704 42944 15784
rect 42944 15704 43024 15784
rect 43024 15704 43104 15784
rect 43104 15704 43184 15784
rect 43184 15704 43264 15784
rect 43264 15704 43344 15784
rect 43344 15704 43424 15784
rect 43424 15704 43504 15784
rect 43504 15704 43584 15784
rect 43584 15704 43664 15784
rect 43664 15704 43744 15784
rect 43744 15704 43824 15784
rect 43824 15704 43904 15784
rect 43904 15704 43984 15784
rect 43984 15704 44064 15784
rect 44064 15704 44144 15784
rect 44144 15704 44224 15784
rect 44224 15704 44304 15784
rect 44304 15704 44384 15784
rect 44384 15704 44464 15784
rect 44464 15704 44544 15784
rect 44544 15704 44624 15784
rect 44624 15704 44704 15784
rect 44704 15704 44784 15784
rect 44784 15704 44864 15784
rect 44864 15704 44944 15784
rect 44944 15704 45024 15784
rect 45024 15704 45104 15784
rect 45104 15704 45184 15784
rect 45184 15704 45264 15784
rect 45264 15704 45344 15784
rect 45344 15704 45424 15784
rect 45424 15704 45504 15784
rect 45504 15704 45584 15784
rect 45584 15704 45664 15784
rect 45664 15704 45744 15784
rect 45744 15704 45824 15784
rect 45824 15704 45904 15784
rect 45904 15704 45984 15784
rect 45984 15704 46064 15784
rect 46064 15704 46144 15784
rect 46144 15704 46224 15784
rect 46224 15704 46304 15784
rect 46304 15704 46384 15784
rect 46384 15704 46464 15784
rect 46464 15704 46544 15784
rect 46544 15704 46624 15784
rect 46624 15704 46704 15784
rect 46704 15704 46784 15784
rect 46784 15704 46864 15784
rect 46864 15704 46944 15784
rect 46944 15704 47024 15784
rect 47024 15704 47104 15784
rect 47104 15704 47184 15784
rect 47184 15704 47264 15784
rect 47264 15704 47344 15784
rect 47344 15704 47424 15784
rect 47424 15704 47504 15784
rect 47504 15704 47584 15784
rect 47584 15704 47664 15784
rect 47664 15704 47744 15784
rect 47744 15704 47824 15784
rect 47824 15704 47904 15784
rect 47904 15704 47984 15784
rect 47984 15704 48064 15784
rect 48064 15704 48144 15784
rect 48144 15704 48224 15784
rect 48224 15704 48304 15784
rect 48304 15704 48384 15784
rect 48384 15704 48464 15784
rect 48464 15704 48544 15784
rect 48544 15704 48624 15784
rect 48624 15704 48704 15784
rect 48704 15704 48784 15784
rect 48784 15704 48864 15784
rect 48864 15704 48944 15784
rect 48944 15704 49024 15784
rect 49024 15704 49104 15784
rect 49104 15704 49184 15784
rect 49184 15704 49264 15784
rect 49264 15704 49344 15784
rect 49344 15704 49424 15784
rect 49424 15704 49504 15784
rect 49504 15704 49584 15784
rect 49584 15704 49664 15784
rect 49664 15704 49744 15784
rect 49744 15704 49824 15784
rect 49824 15704 49904 15784
rect 49904 15704 49984 15784
rect 49984 15704 50064 15784
rect 50064 15704 50144 15784
rect 50144 15704 50224 15784
rect 50224 15704 50304 15784
rect 32 148 112 228
rect 32 228 112 308
rect 32 308 112 388
rect 32 388 112 468
rect 32 468 112 548
rect 32 548 112 628
rect 32 628 112 708
rect 32 708 112 788
rect 32 788 112 868
rect 32 868 112 948
rect 32 948 112 1028
rect 32 1028 112 1108
rect 32 1108 112 1188
rect 32 1188 112 1268
rect 32 1268 112 1348
rect 32 1348 112 1428
rect 32 1428 112 1508
rect 32 1508 112 1588
rect 32 1588 112 1668
rect 32 1668 112 1748
rect 32 1748 112 1828
rect 32 1828 112 1908
rect 32 1908 112 1988
rect 32 1988 112 2068
rect 32 2068 112 2148
rect 32 2148 112 2228
rect 32 2228 112 2308
rect 32 2308 112 2388
rect 32 2388 112 2468
rect 32 2468 112 2548
rect 32 2548 112 2628
rect 32 2628 112 2708
rect 32 2708 112 2788
rect 32 2788 112 2868
rect 32 2868 112 2948
rect 32 2948 112 3028
rect 32 3028 112 3108
rect 32 3108 112 3188
rect 32 3188 112 3268
rect 32 3268 112 3348
rect 32 3348 112 3428
rect 32 3428 112 3508
rect 32 3508 112 3588
rect 32 3588 112 3668
rect 32 3668 112 3748
rect 32 3748 112 3828
rect 32 3828 112 3908
rect 32 3908 112 3988
rect 32 3988 112 4068
rect 32 4068 112 4148
rect 32 4148 112 4228
rect 32 4228 112 4308
rect 32 4308 112 4388
rect 32 4388 112 4468
rect 32 4468 112 4548
rect 32 4548 112 4628
rect 32 4628 112 4708
rect 32 4708 112 4788
rect 32 4788 112 4868
rect 32 4868 112 4948
rect 32 4948 112 5028
rect 32 5028 112 5108
rect 32 5108 112 5188
rect 32 5188 112 5268
rect 32 5268 112 5348
rect 32 5348 112 5428
rect 32 5428 112 5508
rect 32 5508 112 5588
rect 32 5588 112 5668
rect 32 5668 112 5748
rect 32 5748 112 5828
rect 32 5828 112 5908
rect 32 5908 112 5988
rect 32 5988 112 6068
rect 32 6068 112 6148
rect 32 6148 112 6228
rect 32 6228 112 6308
rect 32 6308 112 6388
rect 32 6388 112 6468
rect 32 6468 112 6548
rect 32 6548 112 6628
rect 32 6628 112 6708
rect 32 6708 112 6788
rect 32 6788 112 6868
rect 32 6868 112 6948
rect 32 6948 112 7028
rect 32 7028 112 7108
rect 32 7108 112 7188
rect 32 7188 112 7268
rect 32 7268 112 7348
rect 32 7348 112 7428
rect 32 7428 112 7508
rect 32 7508 112 7588
rect 32 7588 112 7668
rect 32 7668 112 7748
rect 32 7748 112 7828
rect 32 7828 112 7908
rect 32 7908 112 7988
rect 32 7988 112 8068
rect 32 8068 112 8148
rect 32 8148 112 8228
rect 32 8228 112 8308
rect 32 8308 112 8388
rect 32 8388 112 8468
rect 32 8468 112 8548
rect 32 8548 112 8628
rect 32 8628 112 8708
rect 32 8708 112 8788
rect 32 8788 112 8868
rect 32 8868 112 8948
rect 32 8948 112 9028
rect 32 9028 112 9108
rect 32 9108 112 9188
rect 32 9188 112 9268
rect 32 9268 112 9348
rect 32 9348 112 9428
rect 32 9428 112 9508
rect 32 9508 112 9588
rect 32 9588 112 9668
rect 32 9668 112 9748
rect 32 9748 112 9828
rect 32 9828 112 9908
rect 32 9908 112 9988
rect 32 9988 112 10068
rect 32 10068 112 10148
rect 32 10148 112 10228
rect 32 10228 112 10308
rect 32 10308 112 10388
rect 32 10388 112 10468
rect 32 10468 112 10548
rect 32 10548 112 10628
rect 32 10628 112 10708
rect 32 10708 112 10788
rect 32 10788 112 10868
rect 32 10868 112 10948
rect 32 10948 112 11028
rect 32 11028 112 11108
rect 32 11108 112 11188
rect 32 11188 112 11268
rect 32 11268 112 11348
rect 32 11348 112 11428
rect 32 11428 112 11508
rect 32 11508 112 11588
rect 32 11588 112 11668
rect 32 11668 112 11748
rect 32 11748 112 11828
rect 32 11828 112 11908
rect 32 11908 112 11988
rect 32 11988 112 12068
rect 32 12068 112 12148
rect 32 12148 112 12228
rect 32 12228 112 12308
rect 32 12308 112 12388
rect 32 12388 112 12468
rect 32 12468 112 12548
rect 32 12548 112 12628
rect 32 12628 112 12708
rect 32 12708 112 12788
rect 32 12788 112 12868
rect 32 12868 112 12948
rect 32 12948 112 13028
rect 32 13028 112 13108
rect 32 13108 112 13188
rect 32 13188 112 13268
rect 32 13268 112 13348
rect 32 13348 112 13428
rect 32 13428 112 13508
rect 32 13508 112 13588
rect 32 13588 112 13668
rect 32 13668 112 13748
rect 32 13748 112 13828
rect 32 13828 112 13908
rect 32 13908 112 13988
rect 32 13988 112 14068
rect 32 14068 112 14148
rect 32 14148 112 14228
rect 32 14228 112 14308
rect 32 14308 112 14388
rect 32 14388 112 14468
rect 32 14468 112 14548
rect 32 14548 112 14628
rect 32 14628 112 14708
rect 32 14708 112 14788
rect 32 14788 112 14868
rect 32 14868 112 14948
rect 32 14948 112 15028
rect 32 15028 112 15108
rect 32 15108 112 15188
rect 32 15188 112 15268
rect 32 15268 112 15348
rect 32 15348 112 15428
rect 32 15428 112 15508
rect 32 15508 112 15588
rect 32 15588 112 15668
rect 50336 148 50416 228
rect 50336 228 50416 308
rect 50336 308 50416 388
rect 50336 388 50416 468
rect 50336 468 50416 548
rect 50336 548 50416 628
rect 50336 628 50416 708
rect 50336 708 50416 788
rect 50336 788 50416 868
rect 50336 868 50416 948
rect 50336 948 50416 1028
rect 50336 1028 50416 1108
rect 50336 1108 50416 1188
rect 50336 1188 50416 1268
rect 50336 1268 50416 1348
rect 50336 1348 50416 1428
rect 50336 1428 50416 1508
rect 50336 1508 50416 1588
rect 50336 1588 50416 1668
rect 50336 1668 50416 1748
rect 50336 1748 50416 1828
rect 50336 1828 50416 1908
rect 50336 1908 50416 1988
rect 50336 1988 50416 2068
rect 50336 2068 50416 2148
rect 50336 2148 50416 2228
rect 50336 2228 50416 2308
rect 50336 2308 50416 2388
rect 50336 2388 50416 2468
rect 50336 2468 50416 2548
rect 50336 2548 50416 2628
rect 50336 2628 50416 2708
rect 50336 2708 50416 2788
rect 50336 2788 50416 2868
rect 50336 2868 50416 2948
rect 50336 2948 50416 3028
rect 50336 3028 50416 3108
rect 50336 3108 50416 3188
rect 50336 3188 50416 3268
rect 50336 3268 50416 3348
rect 50336 3348 50416 3428
rect 50336 3428 50416 3508
rect 50336 3508 50416 3588
rect 50336 3588 50416 3668
rect 50336 3668 50416 3748
rect 50336 3748 50416 3828
rect 50336 3828 50416 3908
rect 50336 3908 50416 3988
rect 50336 3988 50416 4068
rect 50336 4068 50416 4148
rect 50336 4148 50416 4228
rect 50336 4228 50416 4308
rect 50336 4308 50416 4388
rect 50336 4388 50416 4468
rect 50336 4468 50416 4548
rect 50336 4548 50416 4628
rect 50336 4628 50416 4708
rect 50336 4708 50416 4788
rect 50336 4788 50416 4868
rect 50336 4868 50416 4948
rect 50336 4948 50416 5028
rect 50336 5028 50416 5108
rect 50336 5108 50416 5188
rect 50336 5188 50416 5268
rect 50336 5268 50416 5348
rect 50336 5348 50416 5428
rect 50336 5428 50416 5508
rect 50336 5508 50416 5588
rect 50336 5588 50416 5668
rect 50336 5668 50416 5748
rect 50336 5748 50416 5828
rect 50336 5828 50416 5908
rect 50336 5908 50416 5988
rect 50336 5988 50416 6068
rect 50336 6068 50416 6148
rect 50336 6148 50416 6228
rect 50336 6228 50416 6308
rect 50336 6308 50416 6388
rect 50336 6388 50416 6468
rect 50336 6468 50416 6548
rect 50336 6548 50416 6628
rect 50336 6628 50416 6708
rect 50336 6708 50416 6788
rect 50336 6788 50416 6868
rect 50336 6868 50416 6948
rect 50336 6948 50416 7028
rect 50336 7028 50416 7108
rect 50336 7108 50416 7188
rect 50336 7188 50416 7268
rect 50336 7268 50416 7348
rect 50336 7348 50416 7428
rect 50336 7428 50416 7508
rect 50336 7508 50416 7588
rect 50336 7588 50416 7668
rect 50336 7668 50416 7748
rect 50336 7748 50416 7828
rect 50336 7828 50416 7908
rect 50336 7908 50416 7988
rect 50336 7988 50416 8068
rect 50336 8068 50416 8148
rect 50336 8148 50416 8228
rect 50336 8228 50416 8308
rect 50336 8308 50416 8388
rect 50336 8388 50416 8468
rect 50336 8468 50416 8548
rect 50336 8548 50416 8628
rect 50336 8628 50416 8708
rect 50336 8708 50416 8788
rect 50336 8788 50416 8868
rect 50336 8868 50416 8948
rect 50336 8948 50416 9028
rect 50336 9028 50416 9108
rect 50336 9108 50416 9188
rect 50336 9188 50416 9268
rect 50336 9268 50416 9348
rect 50336 9348 50416 9428
rect 50336 9428 50416 9508
rect 50336 9508 50416 9588
rect 50336 9588 50416 9668
rect 50336 9668 50416 9748
rect 50336 9748 50416 9828
rect 50336 9828 50416 9908
rect 50336 9908 50416 9988
rect 50336 9988 50416 10068
rect 50336 10068 50416 10148
rect 50336 10148 50416 10228
rect 50336 10228 50416 10308
rect 50336 10308 50416 10388
rect 50336 10388 50416 10468
rect 50336 10468 50416 10548
rect 50336 10548 50416 10628
rect 50336 10628 50416 10708
rect 50336 10708 50416 10788
rect 50336 10788 50416 10868
rect 50336 10868 50416 10948
rect 50336 10948 50416 11028
rect 50336 11028 50416 11108
rect 50336 11108 50416 11188
rect 50336 11188 50416 11268
rect 50336 11268 50416 11348
rect 50336 11348 50416 11428
rect 50336 11428 50416 11508
rect 50336 11508 50416 11588
rect 50336 11588 50416 11668
rect 50336 11668 50416 11748
rect 50336 11748 50416 11828
rect 50336 11828 50416 11908
rect 50336 11908 50416 11988
rect 50336 11988 50416 12068
rect 50336 12068 50416 12148
rect 50336 12148 50416 12228
rect 50336 12228 50416 12308
rect 50336 12308 50416 12388
rect 50336 12388 50416 12468
rect 50336 12468 50416 12548
rect 50336 12548 50416 12628
rect 50336 12628 50416 12708
rect 50336 12708 50416 12788
rect 50336 12788 50416 12868
rect 50336 12868 50416 12948
rect 50336 12948 50416 13028
rect 50336 13028 50416 13108
rect 50336 13108 50416 13188
rect 50336 13188 50416 13268
rect 50336 13268 50416 13348
rect 50336 13348 50416 13428
rect 50336 13428 50416 13508
rect 50336 13508 50416 13588
rect 50336 13588 50416 13668
rect 50336 13668 50416 13748
rect 50336 13748 50416 13828
rect 50336 13828 50416 13908
rect 50336 13908 50416 13988
rect 50336 13988 50416 14068
rect 50336 14068 50416 14148
rect 50336 14148 50416 14228
rect 50336 14228 50416 14308
rect 50336 14308 50416 14388
rect 50336 14388 50416 14468
rect 50336 14468 50416 14548
rect 50336 14548 50416 14628
rect 50336 14628 50416 14708
rect 50336 14708 50416 14788
rect 50336 14788 50416 14868
rect 50336 14868 50416 14948
rect 50336 14948 50416 15028
rect 50336 15028 50416 15108
rect 50336 15108 50416 15188
rect 50336 15188 50416 15268
rect 50336 15268 50416 15348
rect 50336 15348 50416 15428
rect 50336 15428 50416 15508
rect 50336 15508 50416 15588
rect 50336 15588 50416 15668
<< ptap >>
rect 0 0 50448 144
rect 0 15672 50448 15816
rect 0 0 144 15816
rect 50304 0 50448 15816
use RPLYBS_PCM XA010
transform 1 0 924 0 1 1364
box 924 1364 2868 12452
use RPLYBS_PCM XA011
transform 1 0 2868 0 1 1364
box 2868 1364 4812 12452
use RPLYBS_PCM XA012
transform 1 0 4812 0 1 1364
box 4812 1364 6756 12452
use RPLYBS_PCM XA013
transform 1 0 6756 0 1 1364
box 6756 1364 8700 12452
use RPLYBS_PCM XB020
transform 1 0 8700 0 1 1364
box 8700 1364 10644 12452
use RPLYBS_PCM XC030
transform 1 0 10644 0 1 1364
box 10644 1364 12588 12452
use RPLYBS_PCM XC031
transform 1 0 12588 0 1 1364
box 12588 1364 14532 12452
use RPLYBS_PCM XC032
transform 1 0 14532 0 1 1364
box 14532 1364 16476 12452
use RPLYBS_PCM XC033
transform 1 0 16476 0 1 1364
box 16476 1364 18420 12452
use RPLYBS_PCM XD040
transform 1 0 18420 0 1 1364
box 18420 1364 20364 12452
use RPLYBS_PCM XD041
transform 1 0 20364 0 1 1364
box 20364 1364 22308 12452
use RPLYBS_PCM XD042
transform 1 0 22308 0 1 1364
box 22308 1364 24252 12452
use RPLYBS_PCM XD043
transform 1 0 24252 0 1 1364
box 24252 1364 26196 12452
use RPLYBS_PCM XB02a0
transform 1 0 26196 0 1 1364
box 26196 1364 28140 12452
use RPLYBS_PCM XF060
transform 1 0 28140 0 1 1364
box 28140 1364 30084 12452
use RPLYBS_PCM XF061
transform 1 0 30084 0 1 1364
box 30084 1364 32028 12452
use RPLYBS_PCM XF062
transform 1 0 32028 0 1 1364
box 32028 1364 33972 12452
use RPLYBS_PCM XF063
transform 1 0 33972 0 1 1364
box 33972 1364 35916 12452
use RPLYBS_PCM XG05a
transform 1 0 35916 0 1 1364
box 35916 1364 37860 12452
use RPLYBS_PCM XG05
transform 1 0 37860 0 1 1364
box 37860 1364 39804 12452
use RPLYBS_PCM XG07
transform 1 0 39804 0 1 1364
box 39804 1364 41748 12452
use RPLYBS_PCM XH08
transform 1 0 41748 0 1 1364
box 41748 1364 43692 12452
use RPLYBS_PCM XI09
transform 1 0 43692 0 1 1364
box 43692 1364 45636 12452
use RPLYBS_PCM XJ10
transform 1 0 45636 0 1 1364
box 45636 1364 47580 12452
use RPLYBS_PCM XK11
transform 1 0 47580 0 1 1364
box 47580 1364 49524 12452
use RPLYBS_cut_M1M4_2x1 
transform 1 0 2336 0 1 5808
box 2336 5808 2536 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 2336 0 1 924
box 2336 924 2536 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 4280 0 1 5808
box 4280 5808 4480 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 4280 0 1 924
box 4280 924 4480 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 6224 0 1 5808
box 6224 5808 6424 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 6224 0 1 924
box 6224 924 6424 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 8168 0 1 5808
box 8168 5808 8368 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 8168 0 1 924
box 8168 924 8368 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 10112 0 1 5808
box 10112 5808 10312 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 10112 0 1 924
box 10112 924 10312 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 12056 0 1 5808
box 12056 5808 12256 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 12056 0 1 924
box 12056 924 12256 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 14000 0 1 5808
box 14000 5808 14200 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 14000 0 1 924
box 14000 924 14200 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 15944 0 1 5808
box 15944 5808 16144 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 15944 0 1 924
box 15944 924 16144 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 17888 0 1 5808
box 17888 5808 18088 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 17888 0 1 924
box 17888 924 18088 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 19832 0 1 5808
box 19832 5808 20032 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 19832 0 1 924
box 19832 924 20032 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 21776 0 1 5808
box 21776 5808 21976 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 21776 0 1 924
box 21776 924 21976 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 23720 0 1 5808
box 23720 5808 23920 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 23720 0 1 924
box 23720 924 23920 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 25664 0 1 5808
box 25664 5808 25864 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 25664 0 1 924
box 25664 924 25864 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 27608 0 1 5808
box 27608 5808 27808 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 27608 0 1 924
box 27608 924 27808 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 29552 0 1 5808
box 29552 5808 29752 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 29552 0 1 924
box 29552 924 29752 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 31496 0 1 5808
box 31496 5808 31696 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 31496 0 1 924
box 31496 924 31696 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 33440 0 1 5808
box 33440 5808 33640 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 33440 0 1 924
box 33440 924 33640 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 35384 0 1 5808
box 35384 5808 35584 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 35384 0 1 924
box 35384 924 35584 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 36384 0 1 8800
box 36384 8800 36584 8876
use RPLYBS_cut_M3M4_2x1 
transform 1 0 36384 0 1 924
box 36384 924 36584 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 37328 0 1 5808
box 37328 5808 37528 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 37328 0 1 924
box 37328 924 37528 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 39272 0 1 5808
box 39272 5808 39472 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 39272 0 1 924
box 39272 924 39472 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 41216 0 1 5808
box 41216 5808 41416 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 41216 0 1 924
box 41216 924 41416 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 43160 0 1 5808
box 43160 5808 43360 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 43160 0 1 924
box 43160 924 43360 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 45104 0 1 5808
box 45104 5808 45304 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 45104 0 1 924
box 45104 924 45304 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 47048 0 1 5808
box 47048 5808 47248 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 47048 0 1 924
box 47048 924 47248 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 48992 0 1 5808
box 48992 5808 49192 5884
use RPLYBS_cut_M3M4_2x1 
transform 1 0 48992 0 1 924
box 48992 924 49192 1000
use RPLYBS_cut_M1M2_2x1 
transform 1 0 2344 0 1 8976
box 2344 8976 2528 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 2336 0 1 12740
box 2336 12740 2536 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 4288 0 1 8976
box 4288 8976 4472 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 4280 0 1 12740
box 4280 12740 4480 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 6232 0 1 8976
box 6232 8976 6416 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 6224 0 1 12740
box 6224 12740 6424 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 8176 0 1 8976
box 8176 8976 8360 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 8168 0 1 12740
box 8168 12740 8368 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 10120 0 1 8976
box 10120 8976 10304 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 10112 0 1 12740
box 10112 12740 10312 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 12064 0 1 8976
box 12064 8976 12248 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 12056 0 1 12740
box 12056 12740 12256 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 14008 0 1 8976
box 14008 8976 14192 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 14000 0 1 12740
box 14000 12740 14200 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 15952 0 1 8976
box 15952 8976 16136 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 15944 0 1 12740
box 15944 12740 16144 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 17896 0 1 8976
box 17896 8976 18080 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 17888 0 1 12740
box 17888 12740 18088 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 19840 0 1 8976
box 19840 8976 20024 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 19832 0 1 12740
box 19832 12740 20032 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 21784 0 1 8976
box 21784 8976 21968 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 21776 0 1 12740
box 21776 12740 21976 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 23728 0 1 8976
box 23728 8976 23912 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 23720 0 1 12740
box 23720 12740 23920 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 25672 0 1 8976
box 25672 8976 25856 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 25664 0 1 12740
box 25664 12740 25864 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 27616 0 1 8976
box 27616 8976 27800 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 27608 0 1 12740
box 27608 12740 27808 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 29560 0 1 8976
box 29560 8976 29744 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 29552 0 1 12740
box 29552 12740 29752 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 31504 0 1 8976
box 31504 8976 31688 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 31496 0 1 12740
box 31496 12740 31696 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 33448 0 1 8976
box 33448 8976 33632 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 33440 0 1 12740
box 33440 12740 33640 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 35392 0 1 8976
box 35392 8976 35576 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 35384 0 1 12740
box 35384 12740 35584 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 37336 0 1 8976
box 37336 8976 37520 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 37328 0 1 12740
box 37328 12740 37528 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 39280 0 1 8976
box 39280 8976 39464 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 39272 0 1 12740
box 39272 12740 39472 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 41224 0 1 8976
box 41224 8976 41408 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 41216 0 1 12740
box 41216 12740 41416 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 43168 0 1 8976
box 43168 8976 43352 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 43160 0 1 12740
box 43160 12740 43360 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 45112 0 1 8976
box 45112 8976 45296 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 45104 0 1 12740
box 45104 12740 45304 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 47056 0 1 8976
box 47056 8976 47240 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 47048 0 1 12740
box 47048 12740 47248 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 49000 0 1 8976
box 49000 8976 49184 9044
use RPLYBS_cut_M2M3_2x1 
transform 1 0 48992 0 1 12740
box 48992 12740 49192 12816
use RPLYBS_cut_M1M2_2x1 
transform 1 0 1392 0 1 8800
box 1392 8800 1576 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 1384 0 1 13768
box 1384 13768 1584 13844
use RPLYBS_cut_M1M2_2x1 
transform 1 0 3336 0 1 8800
box 3336 8800 3520 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 3328 0 1 13768
box 3328 13768 3528 13844
use RPLYBS_cut_M1M2_2x1 
transform 1 0 5280 0 1 8800
box 5280 8800 5464 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 5272 0 1 13768
box 5272 13768 5472 13844
use RPLYBS_cut_M1M2_2x1 
transform 1 0 7224 0 1 8800
box 7224 8800 7408 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 7216 0 1 13768
box 7216 13768 7416 13844
use RPLYBS_cut_M1M2_2x1 
transform 1 0 11112 0 1 8800
box 11112 8800 11296 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 11104 0 1 13768
box 11104 13768 11304 13844
use RPLYBS_cut_M1M2_2x1 
transform 1 0 13056 0 1 8800
box 13056 8800 13240 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 13048 0 1 13768
box 13048 13768 13248 13844
use RPLYBS_cut_M1M2_2x1 
transform 1 0 15000 0 1 8800
box 15000 8800 15184 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 14992 0 1 13768
box 14992 13768 15192 13844
use RPLYBS_cut_M1M2_2x1 
transform 1 0 16944 0 1 8800
box 16944 8800 17128 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 16936 0 1 13768
box 16936 13768 17136 13844
use RPLYBS_cut_M1M2_2x1 
transform 1 0 18888 0 1 8800
box 18888 8800 19072 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 18880 0 1 13768
box 18880 13768 19080 13844
use RPLYBS_cut_M1M2_2x1 
transform 1 0 20832 0 1 8800
box 20832 8800 21016 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 20824 0 1 13768
box 20824 13768 21024 13844
use RPLYBS_cut_M1M2_2x1 
transform 1 0 22776 0 1 8800
box 22776 8800 22960 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 22768 0 1 13768
box 22768 13768 22968 13844
use RPLYBS_cut_M1M2_2x1 
transform 1 0 24720 0 1 8800
box 24720 8800 24904 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 24712 0 1 13768
box 24712 13768 24912 13844
use RPLYBS_cut_M1M2_2x1 
transform 1 0 28608 0 1 8800
box 28608 8800 28792 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 28600 0 1 13768
box 28600 13768 28800 13844
use RPLYBS_cut_M1M2_2x1 
transform 1 0 30552 0 1 8800
box 30552 8800 30736 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 30544 0 1 13768
box 30544 13768 30744 13844
use RPLYBS_cut_M1M2_2x1 
transform 1 0 32496 0 1 8800
box 32496 8800 32680 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 32488 0 1 13768
box 32488 13768 32688 13844
use RPLYBS_cut_M1M2_2x1 
transform 1 0 34440 0 1 8800
box 34440 8800 34624 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 34432 0 1 13768
box 34432 13768 34632 13844
use RPLYBS_cut_M1M2_2x1 
transform 1 0 9168 0 1 8800
box 9168 8800 9352 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 9160 0 1 14208
box 9160 14208 9360 14284
use RPLYBS_cut_M1M2_2x1 
transform 1 0 26664 0 1 8800
box 26664 8800 26848 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 26656 0 1 14208
box 26656 14208 26856 14284
use RPLYBS_cut_M1M2_2x1 
transform 1 0 40272 0 1 8800
box 40272 8800 40456 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 40264 0 1 14432
box 40264 14432 40464 14508
use RPLYBS_cut_M1M2_2x1 
transform 1 0 42216 0 1 8800
box 42216 8800 42400 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 42208 0 1 14656
box 42208 14656 42408 14732
use RPLYBS_cut_M1M2_2x1 
transform 1 0 44160 0 1 8800
box 44160 8800 44344 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 44152 0 1 14880
box 44152 14880 44352 14956
use RPLYBS_cut_M1M2_2x1 
transform 1 0 46104 0 1 8800
box 46104 8800 46288 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 46096 0 1 15104
box 46096 15104 46296 15180
use RPLYBS_cut_M1M2_2x1 
transform 1 0 48048 0 1 8800
box 48048 8800 48232 8868
use RPLYBS_cut_M2M3_2x1 
transform 1 0 48040 0 1 15328
box 48040 15328 48240 15404
use RPLYBS_cut_M1M3_2x1 
transform 1 0 2328 0 1 2640
box 2328 2640 2528 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 4272 0 1 2640
box 4272 2640 4472 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 6216 0 1 2640
box 6216 2640 6416 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 8160 0 1 2640
box 8160 2640 8360 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 10104 0 1 2640
box 10104 2640 10304 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 12048 0 1 2640
box 12048 2640 12248 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 13992 0 1 2640
box 13992 2640 14192 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 15936 0 1 2640
box 15936 2640 16136 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 17880 0 1 2640
box 17880 2640 18080 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 19824 0 1 2640
box 19824 2640 20024 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 21768 0 1 2640
box 21768 2640 21968 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 23712 0 1 2640
box 23712 2640 23912 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 25656 0 1 2640
box 25656 2640 25856 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 27600 0 1 2640
box 27600 2640 27800 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 29544 0 1 2640
box 29544 2640 29744 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 31488 0 1 2640
box 31488 2640 31688 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 33432 0 1 2640
box 33432 2640 33632 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 35376 0 1 2640
box 35376 2640 35576 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 37320 0 1 2640
box 37320 2640 37520 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 39264 0 1 2640
box 39264 2640 39464 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 41208 0 1 2640
box 41208 2640 41408 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 43152 0 1 2640
box 43152 2640 43352 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 45096 0 1 2640
box 45096 2640 45296 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 47040 0 1 2640
box 47040 2640 47240 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 48984 0 1 2640
box 48984 2640 49184 2716
<< labels >>
flabel m2 s 0 924 48600 1076 0 FreeSans 400 0 0 0 VBP
port 1 nsew
flabel m2 s 0 12740 48600 12892 0 FreeSans 400 0 0 0 VCP
port 2 nsew
flabel locali s 49812 336 50112 13480 0 FreeSans 400 0 0 0 AVDD
port 11 nsew
flabel m2 s 1384 13768 34632 13920 0 FreeSans 400 0 0 0 IBP_A
port 3 nsew
flabel m2 s 9160 14208 26856 14360 0 FreeSans 400 0 0 0 IBP_B
port 4 nsew
flabel m2 s 40264 14432 40464 14584 0 FreeSans 400 0 0 0 IBP_1U<4>
port 6 nsew
flabel m2 s 42208 14656 42408 14808 0 FreeSans 400 0 0 0 IBP_1U<3>
port 7 nsew
flabel m2 s 44152 14880 44352 15032 0 FreeSans 400 0 0 0 IBP_1U<2>
port 8 nsew
flabel m2 s 46096 15104 46296 15256 0 FreeSans 400 0 0 0 IBP_1U<1>
port 9 nsew
flabel m2 s 48040 15328 48240 15480 0 FreeSans 400 0 0 0 IBP_1U<0>
port 10 nsew
flabel locali s 16 16 50432 128 0 FreeSans 400 0 0 0 VSS
port 12 nsew
flabel locali s 38328 8800 39048 8888 0 FreeSans 400 0 0 0 IBP_1U<5>
port 5 nsew
flabel m2 s 0 2640 216 2728 0 FreeSans 400 0 0 0 PWRUP_N
port 13 nsew
<< end >>
