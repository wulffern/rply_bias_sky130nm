magic
tech nmos
magscale 1 2
timestamp 1697061600
<< checkpaint >>
rect 0 0 0 0
use CNRATR_NCH_2C12F0 xncm_a_0 ../CNR_ATR_SKY130NM
transform 1 0 0 0 1 0
box 0 0 0 0
use CNRATR_NCH_2C12F0 xncm_a_1[3:0] ../CNR_ATR_SKY130NM
transform 1 0 1152 0 1 0
box 1152 0 1152 0
use CNRATR_NCH_2C12F0 xncm_a_1[3:0] ../CNR_ATR_SKY130NM
transform 1 0 1152 0 1 2030
box 1152 2030 1152 2030
use CNRATR_NCH_2C12F0 xncm_a_1[3:0] ../CNR_ATR_SKY130NM
transform 1 0 1152 0 1 4060
box 1152 4060 1152 4060
use CNRATR_PCH_8C1F2 xpcm_csc_1 ../CNR_ATR_SKY130NM
transform 1 0 2304 0 1 0
box 2304 0 2304 0
use CNRATR_PCH_8C1F2 xpcm_csc_2 ../CNR_ATR_SKY130NM
transform 1 0 4032 0 1 0
box 4032 0 4032 0
use CNRATR_PCH_8C1F2 xpcm_csc_3 ../CNR_ATR_SKY130NM
transform 1 0 5760 0 1 0
box 5760 0 5760 0
use CNRATR_PCH_8C8F0 xpcm_cs_0[15:0] ../CNR_ATR_SKY130NM
transform 1 0 7488 0 1 0
box 7488 0 7488 0
use CNRATR_PCH_8C8F0 xpcm_cs_0[15:0] ../CNR_ATR_SKY130NM
transform 1 0 7488 0 1 1454
box 7488 1454 7488 1454
use CNRATR_PCH_8C8F0 xpcm_cs_0[15:0] ../CNR_ATR_SKY130NM
transform 1 0 7488 0 1 2908
box 7488 2908 7488 2908
use CNRATR_PCH_8C8F0 xpcm_cs_0[15:0] ../CNR_ATR_SKY130NM
transform 1 0 7488 0 1 4362
box 7488 4362 7488 4362
use CNRATR_PCH_8C8F0 xpcm_cs_0[15:0] ../CNR_ATR_SKY130NM
transform 1 0 7488 0 1 5816
box 7488 5816 7488 5816
use CNRATR_PCH_8C8F0 xpcm_cs_0[15:0] ../CNR_ATR_SKY130NM
transform 1 0 7488 0 1 7270
box 7488 7270 7488 7270
use CNRATR_PCH_8C8F0 xpcm_cs_0[15:0] ../CNR_ATR_SKY130NM
transform 1 0 7488 0 1 8724
box 7488 8724 7488 8724
use CNRATR_PCH_8C8F0 xpcm_cs_0[15:0] ../CNR_ATR_SKY130NM
transform 1 0 7488 0 1 10178
box 7488 10178 7488 10178
use CNRATR_PCH_8C8F0 xpcm_cs_0[15:0] ../CNR_ATR_SKY130NM
transform 1 0 7488 0 1 11632
box 7488 11632 7488 11632
use CNRATR_PCH_8C8F0 xpcm_cs_0[15:0] ../CNR_ATR_SKY130NM
transform 1 0 7488 0 1 13086
box 7488 13086 7488 13086
use CNRATR_PCH_8C8F0 xpcm_cs_0[15:0] ../CNR_ATR_SKY130NM
transform 1 0 7488 0 1 14540
box 7488 14540 7488 14540
use CNRATR_PCH_8C8F0 xpcm_cs_0[15:0] ../CNR_ATR_SKY130NM
transform 1 0 7488 0 1 15994
box 7488 15994 7488 15994
use CNRATR_PCH_8C8F0 xpcm_cs_0[15:0] ../CNR_ATR_SKY130NM
transform 1 0 7488 0 1 17448
box 7488 17448 7488 17448
use CNRATR_PCH_8C8F0 xpcm_cs_0[15:0] ../CNR_ATR_SKY130NM
transform 1 0 7488 0 1 18902
box 7488 18902 7488 18902
use CNRATR_PCH_8C8F0 xpcm_cs_0[15:0] ../CNR_ATR_SKY130NM
transform 1 0 7488 0 1 20356
box 7488 20356 7488 20356
use CNRATR_PCH_8C8F0 xpcm_cs_1[1:0] ../CNR_ATR_SKY130NM
transform 1 0 9216 0 1 0
box 9216 0 9216 0
use CNRATR_PCH_8C8F0 xpcm_cs_2 ../CNR_ATR_SKY130NM
transform 1 0 10944 0 1 0
box 10944 0 10944 0
use CNRATR_PCH_8C8F0 xpcm_cs_3 ../CNR_ATR_SKY130NM
transform 1 0 12672 0 1 0
box 12672 0 12672 0
use CNRATR_PCH_8C8F0 xpcm_cs_5 ../CNR_ATR_SKY130NM
transform 1 0 14400 0 1 0
box 14400 0 14400 0
use CNRATR_PCH_8C8F0 xpcm_cs_6 ../CNR_ATR_SKY130NM
transform 1 0 16128 0 1 0
box 16128 0 16128 0
use CNRATR_PCH_8C8F0 xpcm_cs_4 ../CNR_ATR_SKY130NM
transform 1 0 17856 0 1 0
box 17856 0 17856 0
use CNRATR_PCH_8C1F2 xpcm_csc_0[7:0] ../CNR_ATR_SKY130NM
transform 1 0 19584 0 1 0
box 19584 0 19584 0
use CNRATR_PCH_8C1F2 xpcm_csc_0[7:0] ../CNR_ATR_SKY130NM
transform 1 0 19584 0 1 475
box 19584 475 19584 475
use CNRATR_PCH_8C1F2 xpcm_csc_0[7:0] ../CNR_ATR_SKY130NM
transform 1 0 19584 0 1 950
box 19584 950 19584 950
use CNRATR_PCH_8C1F2 xpcm_csc_0[7:0] ../CNR_ATR_SKY130NM
transform 1 0 19584 0 1 1425
box 19584 1425 19584 1425
use CNRATR_PCH_8C1F2 xpcm_csc_0[7:0] ../CNR_ATR_SKY130NM
transform 1 0 19584 0 1 1900
box 19584 1900 19584 1900
use CNRATR_PCH_8C1F2 xpcm_csc_0[7:0] ../CNR_ATR_SKY130NM
transform 1 0 19584 0 1 2375
box 19584 2375 19584 2375
use CNRATR_PCH_8C1F2 xpcm_csc_0[7:0] ../CNR_ATR_SKY130NM
transform 1 0 19584 0 1 2850
box 19584 2850 19584 2850
use CNRATR_PCH_8C1F2 xpcm_csc_4 ../CNR_ATR_SKY130NM
transform 1 0 21312 0 1 0
box 21312 0 21312 0
use CNRATR_PCH_8C1F2 xpcm_csc_5 ../CNR_ATR_SKY130NM
transform 1 0 23040 0 1 0
box 23040 0 23040 0
use CNRATR_PCH_8C1F2 xpcm_csc_6 ../CNR_ATR_SKY130NM
transform 1 0 24768 0 1 0
box 24768 0 24768 0
use CNRATR_PCH_8C8F0 xpcm_vs_0 ../CNR_ATR_SKY130NM
transform 1 0 26496 0 1 0
box 26496 0 26496 0
use CNRATR_NCH_2C12F0 xncm_a_2[1:0] ../CNR_ATR_SKY130NM
transform 1 0 28224 0 1 0
box 28224 0 28224 0
use CNRATR_PCH_8C2F0 xstartp_b_1 ../CNR_ATR_SKY130NM
transform 1 0 29376 0 1 0
box 29376 0 29376 0
use CNRATR_NCH_2C1F2 xstartn_a_0 ../CNR_ATR_SKY130NM
transform 1 0 31104 0 1 0
box 31104 0 31104 0
use CNRATR_NCH_2C12F0 xncm_a_3 ../CNR_ATR_SKY130NM
transform 1 0 32256 0 1 0
box 32256 0 32256 0
use CNRATR_PCH_8C2F0 xstartp_b_0 ../CNR_ATR_SKY130NM
transform 1 0 33408 0 1 0
box 33408 0 33408 0
use CNRATR_NCH_2C12F0 xstartn_a_1 ../CNR_ATR_SKY130NM
transform 1 0 35136 0 1 0
box 35136 0 35136 0
use CNRATR_PCH_8C8F0 xpcm_vs_1 ../CNR_ATR_SKY130NM
transform 1 0 36288 0 1 0
box 36288 0 36288 0
use CNRATR_PCH_8C8F0 xpcm_vs_2 ../CNR_ATR_SKY130NM
transform 1 0 38016 0 1 0
box 38016 0 38016 0
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 0 0
<< end >>
