*TB_SUN_TR_SKY130NM/TB_NCM

.include ../../../work/xsch/RPLY_BIAS.spice

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD 0   dc 1.8

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------

.ic v(VCP)=0.5

IB1 VBP 0 dc 1u
V2 D2 0 dc 0.5
V3 PWRUP_N 0 dc 0

*Cascode
XM3 VBN PWRUP_N VBP VDD PWRUP_N RPLYBS_PCM
XMP1 VBN VBN VSS VSS RPLYBS_NCHCM
XM23 VCP VBN VSS VSS RPLYBS_NCHCM
XC1 VCP VCP VCP1 VDD RPLYBS_PCHCM
XC2 VCP1 VCP VDD VDD RPLYBS_PCHCM

XM1 VBP VCP VBP VDD PWRUP_N RPLYBS_PCM
XM2 D2 VCP VBP VDD PWRUP_N RPLYBS_PCM


.save i(v2) v(XM1.DCM) v(XM1.DCM) v(VDD)




*----------------------------------------------------------------
* NG0PICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 100p 10n 0
dc IB1 10n 2u 0.1u


write


quit

.endc

.end
