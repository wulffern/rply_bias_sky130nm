magic
tech sky130B
magscale 1 2
timestamp 1675206000
<< checkpaint >>
rect 0 0 1944 3168
<< locali >>
rect 756 924 1248 984
rect 828 308 1248 368
rect 1248 308 1308 984
rect 756 1716 1248 1776
rect 828 1100 1248 1160
rect 1248 1100 1308 1776
rect 756 2508 1248 2568
rect 828 1892 1248 1952
rect 1248 1892 1308 2568
rect 828 2684 1248 2744
rect 1248 2684 1308 2744
rect 1482 484 1542 2948
rect -108 220 108 308
rect 468 2684 1188 2772
rect 1404 484 1620 572
rect 324 132 1188 220
use RPLYBS_PCH X1_S0
transform 1 0 0 0 1 0
box 0 0 1944 792
use RPLYBS_PCH X1_S1
transform 1 0 0 0 1 792
box 0 792 1944 1584
use RPLYBS_PCH X1_S2
transform 1 0 0 0 1 1584
box 0 1584 1944 2376
use RPLYBS_PCH X1_S3
transform 1 0 0 0 1 2376
box 0 2376 1944 3168
<< labels >>
flabel locali s -108 220 108 308 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel locali s 468 2684 1188 2772 0 FreeSans 400 0 0 0 D
port 1 nsew
flabel locali s 1404 484 1620 572 0 FreeSans 400 0 0 0 G
port 2 nsew
flabel locali s 324 132 1188 220 0 FreeSans 400 0 0 0 S
port 3 nsew
<< end >>
