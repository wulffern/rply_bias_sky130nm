magic
tech sky130B
magscale 1 2
timestamp 1675206000
<< checkpaint >>
rect 0 0 48504 22152
<< m2 >>
rect 0 924 46656 1076
rect 924 924 47580 1076
rect 0 19076 46656 19228
rect 924 19076 47580 19228
rect 1384 20104 34632 20256
rect 1384 20104 34632 20256
rect 9160 20544 26856 20696
rect 9160 20544 26856 20696
rect 38320 20768 38520 20920
rect 38320 20768 38520 20920
rect 40264 20992 40464 21144
rect 40264 20992 40464 21144
rect 42208 21216 42408 21368
rect 42208 21216 42408 21368
rect 44152 21440 44352 21592
rect 44152 21440 44352 21592
rect 46096 21664 46296 21816
rect 46096 21664 46296 21816
rect 2436 2640 2608 2716
rect 2608 2640 4380 2716
rect 2608 2640 6324 2716
rect 2608 2640 8268 2716
rect 2608 2640 10212 2716
rect 2608 2640 12156 2716
rect 2608 2640 14100 2716
rect 2608 2640 16044 2716
rect 2608 2640 17988 2716
rect 2608 2640 19932 2716
rect 2608 2640 21876 2716
rect 2608 2640 23820 2716
rect 2608 2640 25764 2716
rect 2608 2640 27708 2716
rect 2608 2640 29652 2716
rect 2608 2640 31596 2716
rect 2608 2640 33540 2716
rect 2608 2640 35484 2716
rect 2608 2640 37428 2716
rect 2608 2640 39372 2716
rect 2608 2640 41316 2716
rect 2608 2640 43260 2716
rect 2608 2640 45204 2716
rect 2608 2640 47148 2716
rect 2608 2640 2684 2716
rect 0 2640 216 2728
rect 0 2640 216 2728
rect 2188 2640 2436 2716
rect 108 2640 2188 2716
rect 2188 2640 2264 2716
rect 0 19076 46656 19228
rect 784 19076 24252 19152
rect 784 19076 23328 19152
rect 784 19076 860 19152
rect 0 924 46656 1076
rect 784 924 24252 1000
rect 784 924 23328 1000
rect 784 924 860 1000
<< m3 >>
rect 2398 924 2474 9064
rect 4342 924 4418 9064
rect 6286 924 6362 9064
rect 8230 924 8306 9064
rect 10174 924 10250 9064
rect 12118 924 12194 9064
rect 14062 924 14138 9064
rect 16006 924 16082 9064
rect 17950 924 18026 9064
rect 19894 924 19970 9064
rect 21838 924 21914 9064
rect 23782 924 23858 9064
rect 25726 924 25802 9064
rect 27670 924 27746 9064
rect 29614 924 29690 9064
rect 31558 924 31634 9064
rect 33502 924 33578 9064
rect 35446 924 35522 9064
rect 37390 924 37466 9064
rect 39334 924 39410 9064
rect 41278 924 41354 9064
rect 43222 924 43298 9064
rect 45166 924 45242 9064
rect 47110 924 47186 9064
<< m1 >>
rect 2406 12144 2466 19228
rect 4350 12144 4410 19228
rect 6294 12144 6354 19228
rect 8238 12144 8298 19228
rect 10182 12144 10242 19228
rect 12126 12144 12186 19228
rect 14070 12144 14130 19228
rect 16014 12144 16074 19228
rect 17958 12144 18018 19228
rect 19902 12144 19962 19228
rect 21846 12144 21906 19228
rect 23790 12144 23850 19228
rect 25734 12144 25794 19228
rect 27678 12144 27738 19228
rect 29622 12144 29682 19228
rect 31566 12144 31626 19228
rect 33510 12144 33570 19228
rect 35454 12144 35514 19228
rect 37398 12144 37458 19228
rect 39342 12144 39402 19228
rect 41286 12144 41346 19228
rect 43230 12144 43290 19228
rect 45174 12144 45234 19228
rect 47118 12144 47178 19228
rect 1396 11968 1572 20256
rect 3340 11968 3516 20256
rect 5284 11968 5460 20256
rect 7228 11968 7404 20256
rect 11116 11968 11292 20256
rect 13060 11968 13236 20256
rect 15004 11968 15180 20256
rect 16948 11968 17124 20256
rect 18892 11968 19068 20256
rect 20836 11968 21012 20256
rect 22780 11968 22956 20256
rect 24724 11968 24900 20256
rect 28612 11968 28788 20256
rect 30556 11968 30732 20256
rect 32500 11968 32676 20256
rect 34444 11968 34620 20256
rect 9172 11968 9348 20696
rect 26668 11968 26844 20696
rect 38332 11968 38508 20920
rect 40276 11968 40452 21144
rect 42220 11968 42396 21368
rect 44164 11968 44340 21592
rect 46108 11968 46284 21816
<< locali >>
rect 47868 336 48168 19816
rect 336 336 48168 636
rect 336 19516 48168 19816
rect 336 336 636 19816
rect 47868 336 48168 19816
rect 816 336 1032 1584
rect 816 336 1032 2376
rect 816 336 1032 8712
rect 816 336 1032 11880
rect 816 336 1032 18216
rect 2760 336 2976 1584
rect 2760 336 2976 2376
rect 2760 336 2976 8712
rect 2760 336 2976 11880
rect 2760 336 2976 18216
rect 4704 336 4920 1584
rect 4704 336 4920 2376
rect 4704 336 4920 8712
rect 4704 336 4920 11880
rect 4704 336 4920 18216
rect 6648 336 6864 1584
rect 6648 336 6864 2376
rect 6648 336 6864 8712
rect 6648 336 6864 11880
rect 6648 336 6864 18216
rect 8592 336 8808 1584
rect 8592 336 8808 2376
rect 8592 336 8808 8712
rect 8592 336 8808 11880
rect 8592 336 8808 18216
rect 10536 336 10752 1584
rect 10536 336 10752 2376
rect 10536 336 10752 8712
rect 10536 336 10752 11880
rect 10536 336 10752 18216
rect 12480 336 12696 1584
rect 12480 336 12696 2376
rect 12480 336 12696 8712
rect 12480 336 12696 11880
rect 12480 336 12696 18216
rect 14424 336 14640 1584
rect 14424 336 14640 2376
rect 14424 336 14640 8712
rect 14424 336 14640 11880
rect 14424 336 14640 18216
rect 16368 336 16584 1584
rect 16368 336 16584 2376
rect 16368 336 16584 8712
rect 16368 336 16584 11880
rect 16368 336 16584 18216
rect 18312 336 18528 1584
rect 18312 336 18528 2376
rect 18312 336 18528 8712
rect 18312 336 18528 11880
rect 18312 336 18528 18216
rect 20256 336 20472 1584
rect 20256 336 20472 2376
rect 20256 336 20472 8712
rect 20256 336 20472 11880
rect 20256 336 20472 18216
rect 22200 336 22416 1584
rect 22200 336 22416 2376
rect 22200 336 22416 8712
rect 22200 336 22416 11880
rect 22200 336 22416 18216
rect 24144 336 24360 1584
rect 24144 336 24360 2376
rect 24144 336 24360 8712
rect 24144 336 24360 11880
rect 24144 336 24360 18216
rect 26088 336 26304 1584
rect 26088 336 26304 2376
rect 26088 336 26304 8712
rect 26088 336 26304 11880
rect 26088 336 26304 18216
rect 28032 336 28248 1584
rect 28032 336 28248 2376
rect 28032 336 28248 8712
rect 28032 336 28248 11880
rect 28032 336 28248 18216
rect 29976 336 30192 1584
rect 29976 336 30192 2376
rect 29976 336 30192 8712
rect 29976 336 30192 11880
rect 29976 336 30192 18216
rect 31920 336 32136 1584
rect 31920 336 32136 2376
rect 31920 336 32136 8712
rect 31920 336 32136 11880
rect 31920 336 32136 18216
rect 33864 336 34080 1584
rect 33864 336 34080 2376
rect 33864 336 34080 8712
rect 33864 336 34080 11880
rect 33864 336 34080 18216
rect 35808 336 36024 1584
rect 35808 336 36024 2376
rect 35808 336 36024 8712
rect 35808 336 36024 11880
rect 35808 336 36024 18216
rect 37752 336 37968 1584
rect 37752 336 37968 2376
rect 37752 336 37968 8712
rect 37752 336 37968 11880
rect 37752 336 37968 18216
rect 39696 336 39912 1584
rect 39696 336 39912 2376
rect 39696 336 39912 8712
rect 39696 336 39912 11880
rect 39696 336 39912 18216
rect 41640 336 41856 1584
rect 41640 336 41856 2376
rect 41640 336 41856 8712
rect 41640 336 41856 11880
rect 41640 336 41856 18216
rect 43584 336 43800 1584
rect 43584 336 43800 2376
rect 43584 336 43800 8712
rect 43584 336 43800 11880
rect 43584 336 43800 18216
rect 45528 336 45744 1584
rect 45528 336 45744 2376
rect 45528 336 45744 8712
rect 45528 336 45744 11880
rect 45528 336 45744 18216
rect 16 16 48488 128
rect 128 16 48376 128
rect 128 22024 48376 22136
rect 16 22024 48488 22136
rect 16 128 128 22024
rect 16 16 128 22136
rect 48376 128 48488 22024
rect 48376 16 48488 22136
rect 16 16 48488 128
rect 36384 11968 37104 12056
<< ptapc >>
rect 172 32 252 112
rect 252 32 332 112
rect 332 32 412 112
rect 412 32 492 112
rect 492 32 572 112
rect 572 32 652 112
rect 652 32 732 112
rect 732 32 812 112
rect 812 32 892 112
rect 892 32 972 112
rect 972 32 1052 112
rect 1052 32 1132 112
rect 1132 32 1212 112
rect 1212 32 1292 112
rect 1292 32 1372 112
rect 1372 32 1452 112
rect 1452 32 1532 112
rect 1532 32 1612 112
rect 1612 32 1692 112
rect 1692 32 1772 112
rect 1772 32 1852 112
rect 1852 32 1932 112
rect 1932 32 2012 112
rect 2012 32 2092 112
rect 2092 32 2172 112
rect 2172 32 2252 112
rect 2252 32 2332 112
rect 2332 32 2412 112
rect 2412 32 2492 112
rect 2492 32 2572 112
rect 2572 32 2652 112
rect 2652 32 2732 112
rect 2732 32 2812 112
rect 2812 32 2892 112
rect 2892 32 2972 112
rect 2972 32 3052 112
rect 3052 32 3132 112
rect 3132 32 3212 112
rect 3212 32 3292 112
rect 3292 32 3372 112
rect 3372 32 3452 112
rect 3452 32 3532 112
rect 3532 32 3612 112
rect 3612 32 3692 112
rect 3692 32 3772 112
rect 3772 32 3852 112
rect 3852 32 3932 112
rect 3932 32 4012 112
rect 4012 32 4092 112
rect 4092 32 4172 112
rect 4172 32 4252 112
rect 4252 32 4332 112
rect 4332 32 4412 112
rect 4412 32 4492 112
rect 4492 32 4572 112
rect 4572 32 4652 112
rect 4652 32 4732 112
rect 4732 32 4812 112
rect 4812 32 4892 112
rect 4892 32 4972 112
rect 4972 32 5052 112
rect 5052 32 5132 112
rect 5132 32 5212 112
rect 5212 32 5292 112
rect 5292 32 5372 112
rect 5372 32 5452 112
rect 5452 32 5532 112
rect 5532 32 5612 112
rect 5612 32 5692 112
rect 5692 32 5772 112
rect 5772 32 5852 112
rect 5852 32 5932 112
rect 5932 32 6012 112
rect 6012 32 6092 112
rect 6092 32 6172 112
rect 6172 32 6252 112
rect 6252 32 6332 112
rect 6332 32 6412 112
rect 6412 32 6492 112
rect 6492 32 6572 112
rect 6572 32 6652 112
rect 6652 32 6732 112
rect 6732 32 6812 112
rect 6812 32 6892 112
rect 6892 32 6972 112
rect 6972 32 7052 112
rect 7052 32 7132 112
rect 7132 32 7212 112
rect 7212 32 7292 112
rect 7292 32 7372 112
rect 7372 32 7452 112
rect 7452 32 7532 112
rect 7532 32 7612 112
rect 7612 32 7692 112
rect 7692 32 7772 112
rect 7772 32 7852 112
rect 7852 32 7932 112
rect 7932 32 8012 112
rect 8012 32 8092 112
rect 8092 32 8172 112
rect 8172 32 8252 112
rect 8252 32 8332 112
rect 8332 32 8412 112
rect 8412 32 8492 112
rect 8492 32 8572 112
rect 8572 32 8652 112
rect 8652 32 8732 112
rect 8732 32 8812 112
rect 8812 32 8892 112
rect 8892 32 8972 112
rect 8972 32 9052 112
rect 9052 32 9132 112
rect 9132 32 9212 112
rect 9212 32 9292 112
rect 9292 32 9372 112
rect 9372 32 9452 112
rect 9452 32 9532 112
rect 9532 32 9612 112
rect 9612 32 9692 112
rect 9692 32 9772 112
rect 9772 32 9852 112
rect 9852 32 9932 112
rect 9932 32 10012 112
rect 10012 32 10092 112
rect 10092 32 10172 112
rect 10172 32 10252 112
rect 10252 32 10332 112
rect 10332 32 10412 112
rect 10412 32 10492 112
rect 10492 32 10572 112
rect 10572 32 10652 112
rect 10652 32 10732 112
rect 10732 32 10812 112
rect 10812 32 10892 112
rect 10892 32 10972 112
rect 10972 32 11052 112
rect 11052 32 11132 112
rect 11132 32 11212 112
rect 11212 32 11292 112
rect 11292 32 11372 112
rect 11372 32 11452 112
rect 11452 32 11532 112
rect 11532 32 11612 112
rect 11612 32 11692 112
rect 11692 32 11772 112
rect 11772 32 11852 112
rect 11852 32 11932 112
rect 11932 32 12012 112
rect 12012 32 12092 112
rect 12092 32 12172 112
rect 12172 32 12252 112
rect 12252 32 12332 112
rect 12332 32 12412 112
rect 12412 32 12492 112
rect 12492 32 12572 112
rect 12572 32 12652 112
rect 12652 32 12732 112
rect 12732 32 12812 112
rect 12812 32 12892 112
rect 12892 32 12972 112
rect 12972 32 13052 112
rect 13052 32 13132 112
rect 13132 32 13212 112
rect 13212 32 13292 112
rect 13292 32 13372 112
rect 13372 32 13452 112
rect 13452 32 13532 112
rect 13532 32 13612 112
rect 13612 32 13692 112
rect 13692 32 13772 112
rect 13772 32 13852 112
rect 13852 32 13932 112
rect 13932 32 14012 112
rect 14012 32 14092 112
rect 14092 32 14172 112
rect 14172 32 14252 112
rect 14252 32 14332 112
rect 14332 32 14412 112
rect 14412 32 14492 112
rect 14492 32 14572 112
rect 14572 32 14652 112
rect 14652 32 14732 112
rect 14732 32 14812 112
rect 14812 32 14892 112
rect 14892 32 14972 112
rect 14972 32 15052 112
rect 15052 32 15132 112
rect 15132 32 15212 112
rect 15212 32 15292 112
rect 15292 32 15372 112
rect 15372 32 15452 112
rect 15452 32 15532 112
rect 15532 32 15612 112
rect 15612 32 15692 112
rect 15692 32 15772 112
rect 15772 32 15852 112
rect 15852 32 15932 112
rect 15932 32 16012 112
rect 16012 32 16092 112
rect 16092 32 16172 112
rect 16172 32 16252 112
rect 16252 32 16332 112
rect 16332 32 16412 112
rect 16412 32 16492 112
rect 16492 32 16572 112
rect 16572 32 16652 112
rect 16652 32 16732 112
rect 16732 32 16812 112
rect 16812 32 16892 112
rect 16892 32 16972 112
rect 16972 32 17052 112
rect 17052 32 17132 112
rect 17132 32 17212 112
rect 17212 32 17292 112
rect 17292 32 17372 112
rect 17372 32 17452 112
rect 17452 32 17532 112
rect 17532 32 17612 112
rect 17612 32 17692 112
rect 17692 32 17772 112
rect 17772 32 17852 112
rect 17852 32 17932 112
rect 17932 32 18012 112
rect 18012 32 18092 112
rect 18092 32 18172 112
rect 18172 32 18252 112
rect 18252 32 18332 112
rect 18332 32 18412 112
rect 18412 32 18492 112
rect 18492 32 18572 112
rect 18572 32 18652 112
rect 18652 32 18732 112
rect 18732 32 18812 112
rect 18812 32 18892 112
rect 18892 32 18972 112
rect 18972 32 19052 112
rect 19052 32 19132 112
rect 19132 32 19212 112
rect 19212 32 19292 112
rect 19292 32 19372 112
rect 19372 32 19452 112
rect 19452 32 19532 112
rect 19532 32 19612 112
rect 19612 32 19692 112
rect 19692 32 19772 112
rect 19772 32 19852 112
rect 19852 32 19932 112
rect 19932 32 20012 112
rect 20012 32 20092 112
rect 20092 32 20172 112
rect 20172 32 20252 112
rect 20252 32 20332 112
rect 20332 32 20412 112
rect 20412 32 20492 112
rect 20492 32 20572 112
rect 20572 32 20652 112
rect 20652 32 20732 112
rect 20732 32 20812 112
rect 20812 32 20892 112
rect 20892 32 20972 112
rect 20972 32 21052 112
rect 21052 32 21132 112
rect 21132 32 21212 112
rect 21212 32 21292 112
rect 21292 32 21372 112
rect 21372 32 21452 112
rect 21452 32 21532 112
rect 21532 32 21612 112
rect 21612 32 21692 112
rect 21692 32 21772 112
rect 21772 32 21852 112
rect 21852 32 21932 112
rect 21932 32 22012 112
rect 22012 32 22092 112
rect 22092 32 22172 112
rect 22172 32 22252 112
rect 22252 32 22332 112
rect 22332 32 22412 112
rect 22412 32 22492 112
rect 22492 32 22572 112
rect 22572 32 22652 112
rect 22652 32 22732 112
rect 22732 32 22812 112
rect 22812 32 22892 112
rect 22892 32 22972 112
rect 22972 32 23052 112
rect 23052 32 23132 112
rect 23132 32 23212 112
rect 23212 32 23292 112
rect 23292 32 23372 112
rect 23372 32 23452 112
rect 23452 32 23532 112
rect 23532 32 23612 112
rect 23612 32 23692 112
rect 23692 32 23772 112
rect 23772 32 23852 112
rect 23852 32 23932 112
rect 23932 32 24012 112
rect 24012 32 24092 112
rect 24092 32 24172 112
rect 24172 32 24252 112
rect 24252 32 24332 112
rect 24332 32 24412 112
rect 24412 32 24492 112
rect 24492 32 24572 112
rect 24572 32 24652 112
rect 24652 32 24732 112
rect 24732 32 24812 112
rect 24812 32 24892 112
rect 24892 32 24972 112
rect 24972 32 25052 112
rect 25052 32 25132 112
rect 25132 32 25212 112
rect 25212 32 25292 112
rect 25292 32 25372 112
rect 25372 32 25452 112
rect 25452 32 25532 112
rect 25532 32 25612 112
rect 25612 32 25692 112
rect 25692 32 25772 112
rect 25772 32 25852 112
rect 25852 32 25932 112
rect 25932 32 26012 112
rect 26012 32 26092 112
rect 26092 32 26172 112
rect 26172 32 26252 112
rect 26252 32 26332 112
rect 26332 32 26412 112
rect 26412 32 26492 112
rect 26492 32 26572 112
rect 26572 32 26652 112
rect 26652 32 26732 112
rect 26732 32 26812 112
rect 26812 32 26892 112
rect 26892 32 26972 112
rect 26972 32 27052 112
rect 27052 32 27132 112
rect 27132 32 27212 112
rect 27212 32 27292 112
rect 27292 32 27372 112
rect 27372 32 27452 112
rect 27452 32 27532 112
rect 27532 32 27612 112
rect 27612 32 27692 112
rect 27692 32 27772 112
rect 27772 32 27852 112
rect 27852 32 27932 112
rect 27932 32 28012 112
rect 28012 32 28092 112
rect 28092 32 28172 112
rect 28172 32 28252 112
rect 28252 32 28332 112
rect 28332 32 28412 112
rect 28412 32 28492 112
rect 28492 32 28572 112
rect 28572 32 28652 112
rect 28652 32 28732 112
rect 28732 32 28812 112
rect 28812 32 28892 112
rect 28892 32 28972 112
rect 28972 32 29052 112
rect 29052 32 29132 112
rect 29132 32 29212 112
rect 29212 32 29292 112
rect 29292 32 29372 112
rect 29372 32 29452 112
rect 29452 32 29532 112
rect 29532 32 29612 112
rect 29612 32 29692 112
rect 29692 32 29772 112
rect 29772 32 29852 112
rect 29852 32 29932 112
rect 29932 32 30012 112
rect 30012 32 30092 112
rect 30092 32 30172 112
rect 30172 32 30252 112
rect 30252 32 30332 112
rect 30332 32 30412 112
rect 30412 32 30492 112
rect 30492 32 30572 112
rect 30572 32 30652 112
rect 30652 32 30732 112
rect 30732 32 30812 112
rect 30812 32 30892 112
rect 30892 32 30972 112
rect 30972 32 31052 112
rect 31052 32 31132 112
rect 31132 32 31212 112
rect 31212 32 31292 112
rect 31292 32 31372 112
rect 31372 32 31452 112
rect 31452 32 31532 112
rect 31532 32 31612 112
rect 31612 32 31692 112
rect 31692 32 31772 112
rect 31772 32 31852 112
rect 31852 32 31932 112
rect 31932 32 32012 112
rect 32012 32 32092 112
rect 32092 32 32172 112
rect 32172 32 32252 112
rect 32252 32 32332 112
rect 32332 32 32412 112
rect 32412 32 32492 112
rect 32492 32 32572 112
rect 32572 32 32652 112
rect 32652 32 32732 112
rect 32732 32 32812 112
rect 32812 32 32892 112
rect 32892 32 32972 112
rect 32972 32 33052 112
rect 33052 32 33132 112
rect 33132 32 33212 112
rect 33212 32 33292 112
rect 33292 32 33372 112
rect 33372 32 33452 112
rect 33452 32 33532 112
rect 33532 32 33612 112
rect 33612 32 33692 112
rect 33692 32 33772 112
rect 33772 32 33852 112
rect 33852 32 33932 112
rect 33932 32 34012 112
rect 34012 32 34092 112
rect 34092 32 34172 112
rect 34172 32 34252 112
rect 34252 32 34332 112
rect 34332 32 34412 112
rect 34412 32 34492 112
rect 34492 32 34572 112
rect 34572 32 34652 112
rect 34652 32 34732 112
rect 34732 32 34812 112
rect 34812 32 34892 112
rect 34892 32 34972 112
rect 34972 32 35052 112
rect 35052 32 35132 112
rect 35132 32 35212 112
rect 35212 32 35292 112
rect 35292 32 35372 112
rect 35372 32 35452 112
rect 35452 32 35532 112
rect 35532 32 35612 112
rect 35612 32 35692 112
rect 35692 32 35772 112
rect 35772 32 35852 112
rect 35852 32 35932 112
rect 35932 32 36012 112
rect 36012 32 36092 112
rect 36092 32 36172 112
rect 36172 32 36252 112
rect 36252 32 36332 112
rect 36332 32 36412 112
rect 36412 32 36492 112
rect 36492 32 36572 112
rect 36572 32 36652 112
rect 36652 32 36732 112
rect 36732 32 36812 112
rect 36812 32 36892 112
rect 36892 32 36972 112
rect 36972 32 37052 112
rect 37052 32 37132 112
rect 37132 32 37212 112
rect 37212 32 37292 112
rect 37292 32 37372 112
rect 37372 32 37452 112
rect 37452 32 37532 112
rect 37532 32 37612 112
rect 37612 32 37692 112
rect 37692 32 37772 112
rect 37772 32 37852 112
rect 37852 32 37932 112
rect 37932 32 38012 112
rect 38012 32 38092 112
rect 38092 32 38172 112
rect 38172 32 38252 112
rect 38252 32 38332 112
rect 38332 32 38412 112
rect 38412 32 38492 112
rect 38492 32 38572 112
rect 38572 32 38652 112
rect 38652 32 38732 112
rect 38732 32 38812 112
rect 38812 32 38892 112
rect 38892 32 38972 112
rect 38972 32 39052 112
rect 39052 32 39132 112
rect 39132 32 39212 112
rect 39212 32 39292 112
rect 39292 32 39372 112
rect 39372 32 39452 112
rect 39452 32 39532 112
rect 39532 32 39612 112
rect 39612 32 39692 112
rect 39692 32 39772 112
rect 39772 32 39852 112
rect 39852 32 39932 112
rect 39932 32 40012 112
rect 40012 32 40092 112
rect 40092 32 40172 112
rect 40172 32 40252 112
rect 40252 32 40332 112
rect 40332 32 40412 112
rect 40412 32 40492 112
rect 40492 32 40572 112
rect 40572 32 40652 112
rect 40652 32 40732 112
rect 40732 32 40812 112
rect 40812 32 40892 112
rect 40892 32 40972 112
rect 40972 32 41052 112
rect 41052 32 41132 112
rect 41132 32 41212 112
rect 41212 32 41292 112
rect 41292 32 41372 112
rect 41372 32 41452 112
rect 41452 32 41532 112
rect 41532 32 41612 112
rect 41612 32 41692 112
rect 41692 32 41772 112
rect 41772 32 41852 112
rect 41852 32 41932 112
rect 41932 32 42012 112
rect 42012 32 42092 112
rect 42092 32 42172 112
rect 42172 32 42252 112
rect 42252 32 42332 112
rect 42332 32 42412 112
rect 42412 32 42492 112
rect 42492 32 42572 112
rect 42572 32 42652 112
rect 42652 32 42732 112
rect 42732 32 42812 112
rect 42812 32 42892 112
rect 42892 32 42972 112
rect 42972 32 43052 112
rect 43052 32 43132 112
rect 43132 32 43212 112
rect 43212 32 43292 112
rect 43292 32 43372 112
rect 43372 32 43452 112
rect 43452 32 43532 112
rect 43532 32 43612 112
rect 43612 32 43692 112
rect 43692 32 43772 112
rect 43772 32 43852 112
rect 43852 32 43932 112
rect 43932 32 44012 112
rect 44012 32 44092 112
rect 44092 32 44172 112
rect 44172 32 44252 112
rect 44252 32 44332 112
rect 44332 32 44412 112
rect 44412 32 44492 112
rect 44492 32 44572 112
rect 44572 32 44652 112
rect 44652 32 44732 112
rect 44732 32 44812 112
rect 44812 32 44892 112
rect 44892 32 44972 112
rect 44972 32 45052 112
rect 45052 32 45132 112
rect 45132 32 45212 112
rect 45212 32 45292 112
rect 45292 32 45372 112
rect 45372 32 45452 112
rect 45452 32 45532 112
rect 45532 32 45612 112
rect 45612 32 45692 112
rect 45692 32 45772 112
rect 45772 32 45852 112
rect 45852 32 45932 112
rect 45932 32 46012 112
rect 46012 32 46092 112
rect 46092 32 46172 112
rect 46172 32 46252 112
rect 46252 32 46332 112
rect 46332 32 46412 112
rect 46412 32 46492 112
rect 46492 32 46572 112
rect 46572 32 46652 112
rect 46652 32 46732 112
rect 46732 32 46812 112
rect 46812 32 46892 112
rect 46892 32 46972 112
rect 46972 32 47052 112
rect 47052 32 47132 112
rect 47132 32 47212 112
rect 47212 32 47292 112
rect 47292 32 47372 112
rect 47372 32 47452 112
rect 47452 32 47532 112
rect 47532 32 47612 112
rect 47612 32 47692 112
rect 47692 32 47772 112
rect 47772 32 47852 112
rect 47852 32 47932 112
rect 47932 32 48012 112
rect 48012 32 48092 112
rect 48092 32 48172 112
rect 48172 32 48252 112
rect 48252 32 48332 112
rect 172 22040 252 22120
rect 252 22040 332 22120
rect 332 22040 412 22120
rect 412 22040 492 22120
rect 492 22040 572 22120
rect 572 22040 652 22120
rect 652 22040 732 22120
rect 732 22040 812 22120
rect 812 22040 892 22120
rect 892 22040 972 22120
rect 972 22040 1052 22120
rect 1052 22040 1132 22120
rect 1132 22040 1212 22120
rect 1212 22040 1292 22120
rect 1292 22040 1372 22120
rect 1372 22040 1452 22120
rect 1452 22040 1532 22120
rect 1532 22040 1612 22120
rect 1612 22040 1692 22120
rect 1692 22040 1772 22120
rect 1772 22040 1852 22120
rect 1852 22040 1932 22120
rect 1932 22040 2012 22120
rect 2012 22040 2092 22120
rect 2092 22040 2172 22120
rect 2172 22040 2252 22120
rect 2252 22040 2332 22120
rect 2332 22040 2412 22120
rect 2412 22040 2492 22120
rect 2492 22040 2572 22120
rect 2572 22040 2652 22120
rect 2652 22040 2732 22120
rect 2732 22040 2812 22120
rect 2812 22040 2892 22120
rect 2892 22040 2972 22120
rect 2972 22040 3052 22120
rect 3052 22040 3132 22120
rect 3132 22040 3212 22120
rect 3212 22040 3292 22120
rect 3292 22040 3372 22120
rect 3372 22040 3452 22120
rect 3452 22040 3532 22120
rect 3532 22040 3612 22120
rect 3612 22040 3692 22120
rect 3692 22040 3772 22120
rect 3772 22040 3852 22120
rect 3852 22040 3932 22120
rect 3932 22040 4012 22120
rect 4012 22040 4092 22120
rect 4092 22040 4172 22120
rect 4172 22040 4252 22120
rect 4252 22040 4332 22120
rect 4332 22040 4412 22120
rect 4412 22040 4492 22120
rect 4492 22040 4572 22120
rect 4572 22040 4652 22120
rect 4652 22040 4732 22120
rect 4732 22040 4812 22120
rect 4812 22040 4892 22120
rect 4892 22040 4972 22120
rect 4972 22040 5052 22120
rect 5052 22040 5132 22120
rect 5132 22040 5212 22120
rect 5212 22040 5292 22120
rect 5292 22040 5372 22120
rect 5372 22040 5452 22120
rect 5452 22040 5532 22120
rect 5532 22040 5612 22120
rect 5612 22040 5692 22120
rect 5692 22040 5772 22120
rect 5772 22040 5852 22120
rect 5852 22040 5932 22120
rect 5932 22040 6012 22120
rect 6012 22040 6092 22120
rect 6092 22040 6172 22120
rect 6172 22040 6252 22120
rect 6252 22040 6332 22120
rect 6332 22040 6412 22120
rect 6412 22040 6492 22120
rect 6492 22040 6572 22120
rect 6572 22040 6652 22120
rect 6652 22040 6732 22120
rect 6732 22040 6812 22120
rect 6812 22040 6892 22120
rect 6892 22040 6972 22120
rect 6972 22040 7052 22120
rect 7052 22040 7132 22120
rect 7132 22040 7212 22120
rect 7212 22040 7292 22120
rect 7292 22040 7372 22120
rect 7372 22040 7452 22120
rect 7452 22040 7532 22120
rect 7532 22040 7612 22120
rect 7612 22040 7692 22120
rect 7692 22040 7772 22120
rect 7772 22040 7852 22120
rect 7852 22040 7932 22120
rect 7932 22040 8012 22120
rect 8012 22040 8092 22120
rect 8092 22040 8172 22120
rect 8172 22040 8252 22120
rect 8252 22040 8332 22120
rect 8332 22040 8412 22120
rect 8412 22040 8492 22120
rect 8492 22040 8572 22120
rect 8572 22040 8652 22120
rect 8652 22040 8732 22120
rect 8732 22040 8812 22120
rect 8812 22040 8892 22120
rect 8892 22040 8972 22120
rect 8972 22040 9052 22120
rect 9052 22040 9132 22120
rect 9132 22040 9212 22120
rect 9212 22040 9292 22120
rect 9292 22040 9372 22120
rect 9372 22040 9452 22120
rect 9452 22040 9532 22120
rect 9532 22040 9612 22120
rect 9612 22040 9692 22120
rect 9692 22040 9772 22120
rect 9772 22040 9852 22120
rect 9852 22040 9932 22120
rect 9932 22040 10012 22120
rect 10012 22040 10092 22120
rect 10092 22040 10172 22120
rect 10172 22040 10252 22120
rect 10252 22040 10332 22120
rect 10332 22040 10412 22120
rect 10412 22040 10492 22120
rect 10492 22040 10572 22120
rect 10572 22040 10652 22120
rect 10652 22040 10732 22120
rect 10732 22040 10812 22120
rect 10812 22040 10892 22120
rect 10892 22040 10972 22120
rect 10972 22040 11052 22120
rect 11052 22040 11132 22120
rect 11132 22040 11212 22120
rect 11212 22040 11292 22120
rect 11292 22040 11372 22120
rect 11372 22040 11452 22120
rect 11452 22040 11532 22120
rect 11532 22040 11612 22120
rect 11612 22040 11692 22120
rect 11692 22040 11772 22120
rect 11772 22040 11852 22120
rect 11852 22040 11932 22120
rect 11932 22040 12012 22120
rect 12012 22040 12092 22120
rect 12092 22040 12172 22120
rect 12172 22040 12252 22120
rect 12252 22040 12332 22120
rect 12332 22040 12412 22120
rect 12412 22040 12492 22120
rect 12492 22040 12572 22120
rect 12572 22040 12652 22120
rect 12652 22040 12732 22120
rect 12732 22040 12812 22120
rect 12812 22040 12892 22120
rect 12892 22040 12972 22120
rect 12972 22040 13052 22120
rect 13052 22040 13132 22120
rect 13132 22040 13212 22120
rect 13212 22040 13292 22120
rect 13292 22040 13372 22120
rect 13372 22040 13452 22120
rect 13452 22040 13532 22120
rect 13532 22040 13612 22120
rect 13612 22040 13692 22120
rect 13692 22040 13772 22120
rect 13772 22040 13852 22120
rect 13852 22040 13932 22120
rect 13932 22040 14012 22120
rect 14012 22040 14092 22120
rect 14092 22040 14172 22120
rect 14172 22040 14252 22120
rect 14252 22040 14332 22120
rect 14332 22040 14412 22120
rect 14412 22040 14492 22120
rect 14492 22040 14572 22120
rect 14572 22040 14652 22120
rect 14652 22040 14732 22120
rect 14732 22040 14812 22120
rect 14812 22040 14892 22120
rect 14892 22040 14972 22120
rect 14972 22040 15052 22120
rect 15052 22040 15132 22120
rect 15132 22040 15212 22120
rect 15212 22040 15292 22120
rect 15292 22040 15372 22120
rect 15372 22040 15452 22120
rect 15452 22040 15532 22120
rect 15532 22040 15612 22120
rect 15612 22040 15692 22120
rect 15692 22040 15772 22120
rect 15772 22040 15852 22120
rect 15852 22040 15932 22120
rect 15932 22040 16012 22120
rect 16012 22040 16092 22120
rect 16092 22040 16172 22120
rect 16172 22040 16252 22120
rect 16252 22040 16332 22120
rect 16332 22040 16412 22120
rect 16412 22040 16492 22120
rect 16492 22040 16572 22120
rect 16572 22040 16652 22120
rect 16652 22040 16732 22120
rect 16732 22040 16812 22120
rect 16812 22040 16892 22120
rect 16892 22040 16972 22120
rect 16972 22040 17052 22120
rect 17052 22040 17132 22120
rect 17132 22040 17212 22120
rect 17212 22040 17292 22120
rect 17292 22040 17372 22120
rect 17372 22040 17452 22120
rect 17452 22040 17532 22120
rect 17532 22040 17612 22120
rect 17612 22040 17692 22120
rect 17692 22040 17772 22120
rect 17772 22040 17852 22120
rect 17852 22040 17932 22120
rect 17932 22040 18012 22120
rect 18012 22040 18092 22120
rect 18092 22040 18172 22120
rect 18172 22040 18252 22120
rect 18252 22040 18332 22120
rect 18332 22040 18412 22120
rect 18412 22040 18492 22120
rect 18492 22040 18572 22120
rect 18572 22040 18652 22120
rect 18652 22040 18732 22120
rect 18732 22040 18812 22120
rect 18812 22040 18892 22120
rect 18892 22040 18972 22120
rect 18972 22040 19052 22120
rect 19052 22040 19132 22120
rect 19132 22040 19212 22120
rect 19212 22040 19292 22120
rect 19292 22040 19372 22120
rect 19372 22040 19452 22120
rect 19452 22040 19532 22120
rect 19532 22040 19612 22120
rect 19612 22040 19692 22120
rect 19692 22040 19772 22120
rect 19772 22040 19852 22120
rect 19852 22040 19932 22120
rect 19932 22040 20012 22120
rect 20012 22040 20092 22120
rect 20092 22040 20172 22120
rect 20172 22040 20252 22120
rect 20252 22040 20332 22120
rect 20332 22040 20412 22120
rect 20412 22040 20492 22120
rect 20492 22040 20572 22120
rect 20572 22040 20652 22120
rect 20652 22040 20732 22120
rect 20732 22040 20812 22120
rect 20812 22040 20892 22120
rect 20892 22040 20972 22120
rect 20972 22040 21052 22120
rect 21052 22040 21132 22120
rect 21132 22040 21212 22120
rect 21212 22040 21292 22120
rect 21292 22040 21372 22120
rect 21372 22040 21452 22120
rect 21452 22040 21532 22120
rect 21532 22040 21612 22120
rect 21612 22040 21692 22120
rect 21692 22040 21772 22120
rect 21772 22040 21852 22120
rect 21852 22040 21932 22120
rect 21932 22040 22012 22120
rect 22012 22040 22092 22120
rect 22092 22040 22172 22120
rect 22172 22040 22252 22120
rect 22252 22040 22332 22120
rect 22332 22040 22412 22120
rect 22412 22040 22492 22120
rect 22492 22040 22572 22120
rect 22572 22040 22652 22120
rect 22652 22040 22732 22120
rect 22732 22040 22812 22120
rect 22812 22040 22892 22120
rect 22892 22040 22972 22120
rect 22972 22040 23052 22120
rect 23052 22040 23132 22120
rect 23132 22040 23212 22120
rect 23212 22040 23292 22120
rect 23292 22040 23372 22120
rect 23372 22040 23452 22120
rect 23452 22040 23532 22120
rect 23532 22040 23612 22120
rect 23612 22040 23692 22120
rect 23692 22040 23772 22120
rect 23772 22040 23852 22120
rect 23852 22040 23932 22120
rect 23932 22040 24012 22120
rect 24012 22040 24092 22120
rect 24092 22040 24172 22120
rect 24172 22040 24252 22120
rect 24252 22040 24332 22120
rect 24332 22040 24412 22120
rect 24412 22040 24492 22120
rect 24492 22040 24572 22120
rect 24572 22040 24652 22120
rect 24652 22040 24732 22120
rect 24732 22040 24812 22120
rect 24812 22040 24892 22120
rect 24892 22040 24972 22120
rect 24972 22040 25052 22120
rect 25052 22040 25132 22120
rect 25132 22040 25212 22120
rect 25212 22040 25292 22120
rect 25292 22040 25372 22120
rect 25372 22040 25452 22120
rect 25452 22040 25532 22120
rect 25532 22040 25612 22120
rect 25612 22040 25692 22120
rect 25692 22040 25772 22120
rect 25772 22040 25852 22120
rect 25852 22040 25932 22120
rect 25932 22040 26012 22120
rect 26012 22040 26092 22120
rect 26092 22040 26172 22120
rect 26172 22040 26252 22120
rect 26252 22040 26332 22120
rect 26332 22040 26412 22120
rect 26412 22040 26492 22120
rect 26492 22040 26572 22120
rect 26572 22040 26652 22120
rect 26652 22040 26732 22120
rect 26732 22040 26812 22120
rect 26812 22040 26892 22120
rect 26892 22040 26972 22120
rect 26972 22040 27052 22120
rect 27052 22040 27132 22120
rect 27132 22040 27212 22120
rect 27212 22040 27292 22120
rect 27292 22040 27372 22120
rect 27372 22040 27452 22120
rect 27452 22040 27532 22120
rect 27532 22040 27612 22120
rect 27612 22040 27692 22120
rect 27692 22040 27772 22120
rect 27772 22040 27852 22120
rect 27852 22040 27932 22120
rect 27932 22040 28012 22120
rect 28012 22040 28092 22120
rect 28092 22040 28172 22120
rect 28172 22040 28252 22120
rect 28252 22040 28332 22120
rect 28332 22040 28412 22120
rect 28412 22040 28492 22120
rect 28492 22040 28572 22120
rect 28572 22040 28652 22120
rect 28652 22040 28732 22120
rect 28732 22040 28812 22120
rect 28812 22040 28892 22120
rect 28892 22040 28972 22120
rect 28972 22040 29052 22120
rect 29052 22040 29132 22120
rect 29132 22040 29212 22120
rect 29212 22040 29292 22120
rect 29292 22040 29372 22120
rect 29372 22040 29452 22120
rect 29452 22040 29532 22120
rect 29532 22040 29612 22120
rect 29612 22040 29692 22120
rect 29692 22040 29772 22120
rect 29772 22040 29852 22120
rect 29852 22040 29932 22120
rect 29932 22040 30012 22120
rect 30012 22040 30092 22120
rect 30092 22040 30172 22120
rect 30172 22040 30252 22120
rect 30252 22040 30332 22120
rect 30332 22040 30412 22120
rect 30412 22040 30492 22120
rect 30492 22040 30572 22120
rect 30572 22040 30652 22120
rect 30652 22040 30732 22120
rect 30732 22040 30812 22120
rect 30812 22040 30892 22120
rect 30892 22040 30972 22120
rect 30972 22040 31052 22120
rect 31052 22040 31132 22120
rect 31132 22040 31212 22120
rect 31212 22040 31292 22120
rect 31292 22040 31372 22120
rect 31372 22040 31452 22120
rect 31452 22040 31532 22120
rect 31532 22040 31612 22120
rect 31612 22040 31692 22120
rect 31692 22040 31772 22120
rect 31772 22040 31852 22120
rect 31852 22040 31932 22120
rect 31932 22040 32012 22120
rect 32012 22040 32092 22120
rect 32092 22040 32172 22120
rect 32172 22040 32252 22120
rect 32252 22040 32332 22120
rect 32332 22040 32412 22120
rect 32412 22040 32492 22120
rect 32492 22040 32572 22120
rect 32572 22040 32652 22120
rect 32652 22040 32732 22120
rect 32732 22040 32812 22120
rect 32812 22040 32892 22120
rect 32892 22040 32972 22120
rect 32972 22040 33052 22120
rect 33052 22040 33132 22120
rect 33132 22040 33212 22120
rect 33212 22040 33292 22120
rect 33292 22040 33372 22120
rect 33372 22040 33452 22120
rect 33452 22040 33532 22120
rect 33532 22040 33612 22120
rect 33612 22040 33692 22120
rect 33692 22040 33772 22120
rect 33772 22040 33852 22120
rect 33852 22040 33932 22120
rect 33932 22040 34012 22120
rect 34012 22040 34092 22120
rect 34092 22040 34172 22120
rect 34172 22040 34252 22120
rect 34252 22040 34332 22120
rect 34332 22040 34412 22120
rect 34412 22040 34492 22120
rect 34492 22040 34572 22120
rect 34572 22040 34652 22120
rect 34652 22040 34732 22120
rect 34732 22040 34812 22120
rect 34812 22040 34892 22120
rect 34892 22040 34972 22120
rect 34972 22040 35052 22120
rect 35052 22040 35132 22120
rect 35132 22040 35212 22120
rect 35212 22040 35292 22120
rect 35292 22040 35372 22120
rect 35372 22040 35452 22120
rect 35452 22040 35532 22120
rect 35532 22040 35612 22120
rect 35612 22040 35692 22120
rect 35692 22040 35772 22120
rect 35772 22040 35852 22120
rect 35852 22040 35932 22120
rect 35932 22040 36012 22120
rect 36012 22040 36092 22120
rect 36092 22040 36172 22120
rect 36172 22040 36252 22120
rect 36252 22040 36332 22120
rect 36332 22040 36412 22120
rect 36412 22040 36492 22120
rect 36492 22040 36572 22120
rect 36572 22040 36652 22120
rect 36652 22040 36732 22120
rect 36732 22040 36812 22120
rect 36812 22040 36892 22120
rect 36892 22040 36972 22120
rect 36972 22040 37052 22120
rect 37052 22040 37132 22120
rect 37132 22040 37212 22120
rect 37212 22040 37292 22120
rect 37292 22040 37372 22120
rect 37372 22040 37452 22120
rect 37452 22040 37532 22120
rect 37532 22040 37612 22120
rect 37612 22040 37692 22120
rect 37692 22040 37772 22120
rect 37772 22040 37852 22120
rect 37852 22040 37932 22120
rect 37932 22040 38012 22120
rect 38012 22040 38092 22120
rect 38092 22040 38172 22120
rect 38172 22040 38252 22120
rect 38252 22040 38332 22120
rect 38332 22040 38412 22120
rect 38412 22040 38492 22120
rect 38492 22040 38572 22120
rect 38572 22040 38652 22120
rect 38652 22040 38732 22120
rect 38732 22040 38812 22120
rect 38812 22040 38892 22120
rect 38892 22040 38972 22120
rect 38972 22040 39052 22120
rect 39052 22040 39132 22120
rect 39132 22040 39212 22120
rect 39212 22040 39292 22120
rect 39292 22040 39372 22120
rect 39372 22040 39452 22120
rect 39452 22040 39532 22120
rect 39532 22040 39612 22120
rect 39612 22040 39692 22120
rect 39692 22040 39772 22120
rect 39772 22040 39852 22120
rect 39852 22040 39932 22120
rect 39932 22040 40012 22120
rect 40012 22040 40092 22120
rect 40092 22040 40172 22120
rect 40172 22040 40252 22120
rect 40252 22040 40332 22120
rect 40332 22040 40412 22120
rect 40412 22040 40492 22120
rect 40492 22040 40572 22120
rect 40572 22040 40652 22120
rect 40652 22040 40732 22120
rect 40732 22040 40812 22120
rect 40812 22040 40892 22120
rect 40892 22040 40972 22120
rect 40972 22040 41052 22120
rect 41052 22040 41132 22120
rect 41132 22040 41212 22120
rect 41212 22040 41292 22120
rect 41292 22040 41372 22120
rect 41372 22040 41452 22120
rect 41452 22040 41532 22120
rect 41532 22040 41612 22120
rect 41612 22040 41692 22120
rect 41692 22040 41772 22120
rect 41772 22040 41852 22120
rect 41852 22040 41932 22120
rect 41932 22040 42012 22120
rect 42012 22040 42092 22120
rect 42092 22040 42172 22120
rect 42172 22040 42252 22120
rect 42252 22040 42332 22120
rect 42332 22040 42412 22120
rect 42412 22040 42492 22120
rect 42492 22040 42572 22120
rect 42572 22040 42652 22120
rect 42652 22040 42732 22120
rect 42732 22040 42812 22120
rect 42812 22040 42892 22120
rect 42892 22040 42972 22120
rect 42972 22040 43052 22120
rect 43052 22040 43132 22120
rect 43132 22040 43212 22120
rect 43212 22040 43292 22120
rect 43292 22040 43372 22120
rect 43372 22040 43452 22120
rect 43452 22040 43532 22120
rect 43532 22040 43612 22120
rect 43612 22040 43692 22120
rect 43692 22040 43772 22120
rect 43772 22040 43852 22120
rect 43852 22040 43932 22120
rect 43932 22040 44012 22120
rect 44012 22040 44092 22120
rect 44092 22040 44172 22120
rect 44172 22040 44252 22120
rect 44252 22040 44332 22120
rect 44332 22040 44412 22120
rect 44412 22040 44492 22120
rect 44492 22040 44572 22120
rect 44572 22040 44652 22120
rect 44652 22040 44732 22120
rect 44732 22040 44812 22120
rect 44812 22040 44892 22120
rect 44892 22040 44972 22120
rect 44972 22040 45052 22120
rect 45052 22040 45132 22120
rect 45132 22040 45212 22120
rect 45212 22040 45292 22120
rect 45292 22040 45372 22120
rect 45372 22040 45452 22120
rect 45452 22040 45532 22120
rect 45532 22040 45612 22120
rect 45612 22040 45692 22120
rect 45692 22040 45772 22120
rect 45772 22040 45852 22120
rect 45852 22040 45932 22120
rect 45932 22040 46012 22120
rect 46012 22040 46092 22120
rect 46092 22040 46172 22120
rect 46172 22040 46252 22120
rect 46252 22040 46332 22120
rect 46332 22040 46412 22120
rect 46412 22040 46492 22120
rect 46492 22040 46572 22120
rect 46572 22040 46652 22120
rect 46652 22040 46732 22120
rect 46732 22040 46812 22120
rect 46812 22040 46892 22120
rect 46892 22040 46972 22120
rect 46972 22040 47052 22120
rect 47052 22040 47132 22120
rect 47132 22040 47212 22120
rect 47212 22040 47292 22120
rect 47292 22040 47372 22120
rect 47372 22040 47452 22120
rect 47452 22040 47532 22120
rect 47532 22040 47612 22120
rect 47612 22040 47692 22120
rect 47692 22040 47772 22120
rect 47772 22040 47852 22120
rect 47852 22040 47932 22120
rect 47932 22040 48012 22120
rect 48012 22040 48092 22120
rect 48092 22040 48172 22120
rect 48172 22040 48252 22120
rect 48252 22040 48332 22120
rect 32 156 112 236
rect 32 236 112 316
rect 32 316 112 396
rect 32 396 112 476
rect 32 476 112 556
rect 32 556 112 636
rect 32 636 112 716
rect 32 716 112 796
rect 32 796 112 876
rect 32 876 112 956
rect 32 956 112 1036
rect 32 1036 112 1116
rect 32 1116 112 1196
rect 32 1196 112 1276
rect 32 1276 112 1356
rect 32 1356 112 1436
rect 32 1436 112 1516
rect 32 1516 112 1596
rect 32 1596 112 1676
rect 32 1676 112 1756
rect 32 1756 112 1836
rect 32 1836 112 1916
rect 32 1916 112 1996
rect 32 1996 112 2076
rect 32 2076 112 2156
rect 32 2156 112 2236
rect 32 2236 112 2316
rect 32 2316 112 2396
rect 32 2396 112 2476
rect 32 2476 112 2556
rect 32 2556 112 2636
rect 32 2636 112 2716
rect 32 2716 112 2796
rect 32 2796 112 2876
rect 32 2876 112 2956
rect 32 2956 112 3036
rect 32 3036 112 3116
rect 32 3116 112 3196
rect 32 3196 112 3276
rect 32 3276 112 3356
rect 32 3356 112 3436
rect 32 3436 112 3516
rect 32 3516 112 3596
rect 32 3596 112 3676
rect 32 3676 112 3756
rect 32 3756 112 3836
rect 32 3836 112 3916
rect 32 3916 112 3996
rect 32 3996 112 4076
rect 32 4076 112 4156
rect 32 4156 112 4236
rect 32 4236 112 4316
rect 32 4316 112 4396
rect 32 4396 112 4476
rect 32 4476 112 4556
rect 32 4556 112 4636
rect 32 4636 112 4716
rect 32 4716 112 4796
rect 32 4796 112 4876
rect 32 4876 112 4956
rect 32 4956 112 5036
rect 32 5036 112 5116
rect 32 5116 112 5196
rect 32 5196 112 5276
rect 32 5276 112 5356
rect 32 5356 112 5436
rect 32 5436 112 5516
rect 32 5516 112 5596
rect 32 5596 112 5676
rect 32 5676 112 5756
rect 32 5756 112 5836
rect 32 5836 112 5916
rect 32 5916 112 5996
rect 32 5996 112 6076
rect 32 6076 112 6156
rect 32 6156 112 6236
rect 32 6236 112 6316
rect 32 6316 112 6396
rect 32 6396 112 6476
rect 32 6476 112 6556
rect 32 6556 112 6636
rect 32 6636 112 6716
rect 32 6716 112 6796
rect 32 6796 112 6876
rect 32 6876 112 6956
rect 32 6956 112 7036
rect 32 7036 112 7116
rect 32 7116 112 7196
rect 32 7196 112 7276
rect 32 7276 112 7356
rect 32 7356 112 7436
rect 32 7436 112 7516
rect 32 7516 112 7596
rect 32 7596 112 7676
rect 32 7676 112 7756
rect 32 7756 112 7836
rect 32 7836 112 7916
rect 32 7916 112 7996
rect 32 7996 112 8076
rect 32 8076 112 8156
rect 32 8156 112 8236
rect 32 8236 112 8316
rect 32 8316 112 8396
rect 32 8396 112 8476
rect 32 8476 112 8556
rect 32 8556 112 8636
rect 32 8636 112 8716
rect 32 8716 112 8796
rect 32 8796 112 8876
rect 32 8876 112 8956
rect 32 8956 112 9036
rect 32 9036 112 9116
rect 32 9116 112 9196
rect 32 9196 112 9276
rect 32 9276 112 9356
rect 32 9356 112 9436
rect 32 9436 112 9516
rect 32 9516 112 9596
rect 32 9596 112 9676
rect 32 9676 112 9756
rect 32 9756 112 9836
rect 32 9836 112 9916
rect 32 9916 112 9996
rect 32 9996 112 10076
rect 32 10076 112 10156
rect 32 10156 112 10236
rect 32 10236 112 10316
rect 32 10316 112 10396
rect 32 10396 112 10476
rect 32 10476 112 10556
rect 32 10556 112 10636
rect 32 10636 112 10716
rect 32 10716 112 10796
rect 32 10796 112 10876
rect 32 10876 112 10956
rect 32 10956 112 11036
rect 32 11036 112 11116
rect 32 11116 112 11196
rect 32 11196 112 11276
rect 32 11276 112 11356
rect 32 11356 112 11436
rect 32 11436 112 11516
rect 32 11516 112 11596
rect 32 11596 112 11676
rect 32 11676 112 11756
rect 32 11756 112 11836
rect 32 11836 112 11916
rect 32 11916 112 11996
rect 32 11996 112 12076
rect 32 12076 112 12156
rect 32 12156 112 12236
rect 32 12236 112 12316
rect 32 12316 112 12396
rect 32 12396 112 12476
rect 32 12476 112 12556
rect 32 12556 112 12636
rect 32 12636 112 12716
rect 32 12716 112 12796
rect 32 12796 112 12876
rect 32 12876 112 12956
rect 32 12956 112 13036
rect 32 13036 112 13116
rect 32 13116 112 13196
rect 32 13196 112 13276
rect 32 13276 112 13356
rect 32 13356 112 13436
rect 32 13436 112 13516
rect 32 13516 112 13596
rect 32 13596 112 13676
rect 32 13676 112 13756
rect 32 13756 112 13836
rect 32 13836 112 13916
rect 32 13916 112 13996
rect 32 13996 112 14076
rect 32 14076 112 14156
rect 32 14156 112 14236
rect 32 14236 112 14316
rect 32 14316 112 14396
rect 32 14396 112 14476
rect 32 14476 112 14556
rect 32 14556 112 14636
rect 32 14636 112 14716
rect 32 14716 112 14796
rect 32 14796 112 14876
rect 32 14876 112 14956
rect 32 14956 112 15036
rect 32 15036 112 15116
rect 32 15116 112 15196
rect 32 15196 112 15276
rect 32 15276 112 15356
rect 32 15356 112 15436
rect 32 15436 112 15516
rect 32 15516 112 15596
rect 32 15596 112 15676
rect 32 15676 112 15756
rect 32 15756 112 15836
rect 32 15836 112 15916
rect 32 15916 112 15996
rect 32 15996 112 16076
rect 32 16076 112 16156
rect 32 16156 112 16236
rect 32 16236 112 16316
rect 32 16316 112 16396
rect 32 16396 112 16476
rect 32 16476 112 16556
rect 32 16556 112 16636
rect 32 16636 112 16716
rect 32 16716 112 16796
rect 32 16796 112 16876
rect 32 16876 112 16956
rect 32 16956 112 17036
rect 32 17036 112 17116
rect 32 17116 112 17196
rect 32 17196 112 17276
rect 32 17276 112 17356
rect 32 17356 112 17436
rect 32 17436 112 17516
rect 32 17516 112 17596
rect 32 17596 112 17676
rect 32 17676 112 17756
rect 32 17756 112 17836
rect 32 17836 112 17916
rect 32 17916 112 17996
rect 32 17996 112 18076
rect 32 18076 112 18156
rect 32 18156 112 18236
rect 32 18236 112 18316
rect 32 18316 112 18396
rect 32 18396 112 18476
rect 32 18476 112 18556
rect 32 18556 112 18636
rect 32 18636 112 18716
rect 32 18716 112 18796
rect 32 18796 112 18876
rect 32 18876 112 18956
rect 32 18956 112 19036
rect 32 19036 112 19116
rect 32 19116 112 19196
rect 32 19196 112 19276
rect 32 19276 112 19356
rect 32 19356 112 19436
rect 32 19436 112 19516
rect 32 19516 112 19596
rect 32 19596 112 19676
rect 32 19676 112 19756
rect 32 19756 112 19836
rect 32 19836 112 19916
rect 32 19916 112 19996
rect 32 19996 112 20076
rect 32 20076 112 20156
rect 32 20156 112 20236
rect 32 20236 112 20316
rect 32 20316 112 20396
rect 32 20396 112 20476
rect 32 20476 112 20556
rect 32 20556 112 20636
rect 32 20636 112 20716
rect 32 20716 112 20796
rect 32 20796 112 20876
rect 32 20876 112 20956
rect 32 20956 112 21036
rect 32 21036 112 21116
rect 32 21116 112 21196
rect 32 21196 112 21276
rect 32 21276 112 21356
rect 32 21356 112 21436
rect 32 21436 112 21516
rect 32 21516 112 21596
rect 32 21596 112 21676
rect 32 21676 112 21756
rect 32 21756 112 21836
rect 32 21836 112 21916
rect 32 21916 112 21996
rect 48392 156 48472 236
rect 48392 236 48472 316
rect 48392 316 48472 396
rect 48392 396 48472 476
rect 48392 476 48472 556
rect 48392 556 48472 636
rect 48392 636 48472 716
rect 48392 716 48472 796
rect 48392 796 48472 876
rect 48392 876 48472 956
rect 48392 956 48472 1036
rect 48392 1036 48472 1116
rect 48392 1116 48472 1196
rect 48392 1196 48472 1276
rect 48392 1276 48472 1356
rect 48392 1356 48472 1436
rect 48392 1436 48472 1516
rect 48392 1516 48472 1596
rect 48392 1596 48472 1676
rect 48392 1676 48472 1756
rect 48392 1756 48472 1836
rect 48392 1836 48472 1916
rect 48392 1916 48472 1996
rect 48392 1996 48472 2076
rect 48392 2076 48472 2156
rect 48392 2156 48472 2236
rect 48392 2236 48472 2316
rect 48392 2316 48472 2396
rect 48392 2396 48472 2476
rect 48392 2476 48472 2556
rect 48392 2556 48472 2636
rect 48392 2636 48472 2716
rect 48392 2716 48472 2796
rect 48392 2796 48472 2876
rect 48392 2876 48472 2956
rect 48392 2956 48472 3036
rect 48392 3036 48472 3116
rect 48392 3116 48472 3196
rect 48392 3196 48472 3276
rect 48392 3276 48472 3356
rect 48392 3356 48472 3436
rect 48392 3436 48472 3516
rect 48392 3516 48472 3596
rect 48392 3596 48472 3676
rect 48392 3676 48472 3756
rect 48392 3756 48472 3836
rect 48392 3836 48472 3916
rect 48392 3916 48472 3996
rect 48392 3996 48472 4076
rect 48392 4076 48472 4156
rect 48392 4156 48472 4236
rect 48392 4236 48472 4316
rect 48392 4316 48472 4396
rect 48392 4396 48472 4476
rect 48392 4476 48472 4556
rect 48392 4556 48472 4636
rect 48392 4636 48472 4716
rect 48392 4716 48472 4796
rect 48392 4796 48472 4876
rect 48392 4876 48472 4956
rect 48392 4956 48472 5036
rect 48392 5036 48472 5116
rect 48392 5116 48472 5196
rect 48392 5196 48472 5276
rect 48392 5276 48472 5356
rect 48392 5356 48472 5436
rect 48392 5436 48472 5516
rect 48392 5516 48472 5596
rect 48392 5596 48472 5676
rect 48392 5676 48472 5756
rect 48392 5756 48472 5836
rect 48392 5836 48472 5916
rect 48392 5916 48472 5996
rect 48392 5996 48472 6076
rect 48392 6076 48472 6156
rect 48392 6156 48472 6236
rect 48392 6236 48472 6316
rect 48392 6316 48472 6396
rect 48392 6396 48472 6476
rect 48392 6476 48472 6556
rect 48392 6556 48472 6636
rect 48392 6636 48472 6716
rect 48392 6716 48472 6796
rect 48392 6796 48472 6876
rect 48392 6876 48472 6956
rect 48392 6956 48472 7036
rect 48392 7036 48472 7116
rect 48392 7116 48472 7196
rect 48392 7196 48472 7276
rect 48392 7276 48472 7356
rect 48392 7356 48472 7436
rect 48392 7436 48472 7516
rect 48392 7516 48472 7596
rect 48392 7596 48472 7676
rect 48392 7676 48472 7756
rect 48392 7756 48472 7836
rect 48392 7836 48472 7916
rect 48392 7916 48472 7996
rect 48392 7996 48472 8076
rect 48392 8076 48472 8156
rect 48392 8156 48472 8236
rect 48392 8236 48472 8316
rect 48392 8316 48472 8396
rect 48392 8396 48472 8476
rect 48392 8476 48472 8556
rect 48392 8556 48472 8636
rect 48392 8636 48472 8716
rect 48392 8716 48472 8796
rect 48392 8796 48472 8876
rect 48392 8876 48472 8956
rect 48392 8956 48472 9036
rect 48392 9036 48472 9116
rect 48392 9116 48472 9196
rect 48392 9196 48472 9276
rect 48392 9276 48472 9356
rect 48392 9356 48472 9436
rect 48392 9436 48472 9516
rect 48392 9516 48472 9596
rect 48392 9596 48472 9676
rect 48392 9676 48472 9756
rect 48392 9756 48472 9836
rect 48392 9836 48472 9916
rect 48392 9916 48472 9996
rect 48392 9996 48472 10076
rect 48392 10076 48472 10156
rect 48392 10156 48472 10236
rect 48392 10236 48472 10316
rect 48392 10316 48472 10396
rect 48392 10396 48472 10476
rect 48392 10476 48472 10556
rect 48392 10556 48472 10636
rect 48392 10636 48472 10716
rect 48392 10716 48472 10796
rect 48392 10796 48472 10876
rect 48392 10876 48472 10956
rect 48392 10956 48472 11036
rect 48392 11036 48472 11116
rect 48392 11116 48472 11196
rect 48392 11196 48472 11276
rect 48392 11276 48472 11356
rect 48392 11356 48472 11436
rect 48392 11436 48472 11516
rect 48392 11516 48472 11596
rect 48392 11596 48472 11676
rect 48392 11676 48472 11756
rect 48392 11756 48472 11836
rect 48392 11836 48472 11916
rect 48392 11916 48472 11996
rect 48392 11996 48472 12076
rect 48392 12076 48472 12156
rect 48392 12156 48472 12236
rect 48392 12236 48472 12316
rect 48392 12316 48472 12396
rect 48392 12396 48472 12476
rect 48392 12476 48472 12556
rect 48392 12556 48472 12636
rect 48392 12636 48472 12716
rect 48392 12716 48472 12796
rect 48392 12796 48472 12876
rect 48392 12876 48472 12956
rect 48392 12956 48472 13036
rect 48392 13036 48472 13116
rect 48392 13116 48472 13196
rect 48392 13196 48472 13276
rect 48392 13276 48472 13356
rect 48392 13356 48472 13436
rect 48392 13436 48472 13516
rect 48392 13516 48472 13596
rect 48392 13596 48472 13676
rect 48392 13676 48472 13756
rect 48392 13756 48472 13836
rect 48392 13836 48472 13916
rect 48392 13916 48472 13996
rect 48392 13996 48472 14076
rect 48392 14076 48472 14156
rect 48392 14156 48472 14236
rect 48392 14236 48472 14316
rect 48392 14316 48472 14396
rect 48392 14396 48472 14476
rect 48392 14476 48472 14556
rect 48392 14556 48472 14636
rect 48392 14636 48472 14716
rect 48392 14716 48472 14796
rect 48392 14796 48472 14876
rect 48392 14876 48472 14956
rect 48392 14956 48472 15036
rect 48392 15036 48472 15116
rect 48392 15116 48472 15196
rect 48392 15196 48472 15276
rect 48392 15276 48472 15356
rect 48392 15356 48472 15436
rect 48392 15436 48472 15516
rect 48392 15516 48472 15596
rect 48392 15596 48472 15676
rect 48392 15676 48472 15756
rect 48392 15756 48472 15836
rect 48392 15836 48472 15916
rect 48392 15916 48472 15996
rect 48392 15996 48472 16076
rect 48392 16076 48472 16156
rect 48392 16156 48472 16236
rect 48392 16236 48472 16316
rect 48392 16316 48472 16396
rect 48392 16396 48472 16476
rect 48392 16476 48472 16556
rect 48392 16556 48472 16636
rect 48392 16636 48472 16716
rect 48392 16716 48472 16796
rect 48392 16796 48472 16876
rect 48392 16876 48472 16956
rect 48392 16956 48472 17036
rect 48392 17036 48472 17116
rect 48392 17116 48472 17196
rect 48392 17196 48472 17276
rect 48392 17276 48472 17356
rect 48392 17356 48472 17436
rect 48392 17436 48472 17516
rect 48392 17516 48472 17596
rect 48392 17596 48472 17676
rect 48392 17676 48472 17756
rect 48392 17756 48472 17836
rect 48392 17836 48472 17916
rect 48392 17916 48472 17996
rect 48392 17996 48472 18076
rect 48392 18076 48472 18156
rect 48392 18156 48472 18236
rect 48392 18236 48472 18316
rect 48392 18316 48472 18396
rect 48392 18396 48472 18476
rect 48392 18476 48472 18556
rect 48392 18556 48472 18636
rect 48392 18636 48472 18716
rect 48392 18716 48472 18796
rect 48392 18796 48472 18876
rect 48392 18876 48472 18956
rect 48392 18956 48472 19036
rect 48392 19036 48472 19116
rect 48392 19116 48472 19196
rect 48392 19196 48472 19276
rect 48392 19276 48472 19356
rect 48392 19356 48472 19436
rect 48392 19436 48472 19516
rect 48392 19516 48472 19596
rect 48392 19596 48472 19676
rect 48392 19676 48472 19756
rect 48392 19756 48472 19836
rect 48392 19836 48472 19916
rect 48392 19916 48472 19996
rect 48392 19996 48472 20076
rect 48392 20076 48472 20156
rect 48392 20156 48472 20236
rect 48392 20236 48472 20316
rect 48392 20316 48472 20396
rect 48392 20396 48472 20476
rect 48392 20476 48472 20556
rect 48392 20556 48472 20636
rect 48392 20636 48472 20716
rect 48392 20716 48472 20796
rect 48392 20796 48472 20876
rect 48392 20876 48472 20956
rect 48392 20956 48472 21036
rect 48392 21036 48472 21116
rect 48392 21116 48472 21196
rect 48392 21196 48472 21276
rect 48392 21276 48472 21356
rect 48392 21356 48472 21436
rect 48392 21436 48472 21516
rect 48392 21516 48472 21596
rect 48392 21596 48472 21676
rect 48392 21676 48472 21756
rect 48392 21756 48472 21836
rect 48392 21836 48472 21916
rect 48392 21916 48472 21996
<< ptap >>
rect 0 0 48504 144
rect 0 22008 48504 22152
rect 0 0 144 22152
rect 48360 0 48504 22152
use RPLYBS_PCM XA010
transform 1 0 924 0 1 1364
box 924 1364 2868 18788
use RPLYBS_PCM XA011
transform 1 0 2868 0 1 1364
box 2868 1364 4812 18788
use RPLYBS_PCM XA012
transform 1 0 4812 0 1 1364
box 4812 1364 6756 18788
use RPLYBS_PCM XA013
transform 1 0 6756 0 1 1364
box 6756 1364 8700 18788
use RPLYBS_PCM XB020
transform 1 0 8700 0 1 1364
box 8700 1364 10644 18788
use RPLYBS_PCM XC030
transform 1 0 10644 0 1 1364
box 10644 1364 12588 18788
use RPLYBS_PCM XC031
transform 1 0 12588 0 1 1364
box 12588 1364 14532 18788
use RPLYBS_PCM XC032
transform 1 0 14532 0 1 1364
box 14532 1364 16476 18788
use RPLYBS_PCM XC033
transform 1 0 16476 0 1 1364
box 16476 1364 18420 18788
use RPLYBS_PCM XD040
transform 1 0 18420 0 1 1364
box 18420 1364 20364 18788
use RPLYBS_PCM XD041
transform 1 0 20364 0 1 1364
box 20364 1364 22308 18788
use RPLYBS_PCM XD042
transform 1 0 22308 0 1 1364
box 22308 1364 24252 18788
use RPLYBS_PCM XD043
transform 1 0 24252 0 1 1364
box 24252 1364 26196 18788
use RPLYBS_PCM XE050
transform 1 0 26196 0 1 1364
box 26196 1364 28140 18788
use RPLYBS_PCM XF060
transform 1 0 28140 0 1 1364
box 28140 1364 30084 18788
use RPLYBS_PCM XF061
transform 1 0 30084 0 1 1364
box 30084 1364 32028 18788
use RPLYBS_PCM XF062
transform 1 0 32028 0 1 1364
box 32028 1364 33972 18788
use RPLYBS_PCM XF063
transform 1 0 33972 0 1 1364
box 33972 1364 35916 18788
use RPLYBS_PCM XG05
transform 1 0 35916 0 1 1364
box 35916 1364 37860 18788
use RPLYBS_PCM XG07
transform 1 0 37860 0 1 1364
box 37860 1364 39804 18788
use RPLYBS_PCM XH08
transform 1 0 39804 0 1 1364
box 39804 1364 41748 18788
use RPLYBS_PCM XI09
transform 1 0 41748 0 1 1364
box 41748 1364 43692 18788
use RPLYBS_PCM XJ10
transform 1 0 43692 0 1 1364
box 43692 1364 45636 18788
use RPLYBS_PCM XK11
transform 1 0 45636 0 1 1364
box 45636 1364 47580 18788
use RPLYBS_cut_M1M4_2x1 
transform 1 0 2336 0 1 8976
box 2336 8976 2536 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 2336 0 1 924
box 2336 924 2536 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 4280 0 1 8976
box 4280 8976 4480 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 4280 0 1 924
box 4280 924 4480 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 6224 0 1 8976
box 6224 8976 6424 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 6224 0 1 924
box 6224 924 6424 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 8168 0 1 8976
box 8168 8976 8368 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 8168 0 1 924
box 8168 924 8368 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 10112 0 1 8976
box 10112 8976 10312 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 10112 0 1 924
box 10112 924 10312 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 12056 0 1 8976
box 12056 8976 12256 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 12056 0 1 924
box 12056 924 12256 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 14000 0 1 8976
box 14000 8976 14200 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 14000 0 1 924
box 14000 924 14200 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 15944 0 1 8976
box 15944 8976 16144 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 15944 0 1 924
box 15944 924 16144 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 17888 0 1 8976
box 17888 8976 18088 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 17888 0 1 924
box 17888 924 18088 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 19832 0 1 8976
box 19832 8976 20032 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 19832 0 1 924
box 19832 924 20032 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 21776 0 1 8976
box 21776 8976 21976 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 21776 0 1 924
box 21776 924 21976 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 23720 0 1 8976
box 23720 8976 23920 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 23720 0 1 924
box 23720 924 23920 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 25664 0 1 8976
box 25664 8976 25864 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 25664 0 1 924
box 25664 924 25864 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 27608 0 1 8976
box 27608 8976 27808 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 27608 0 1 924
box 27608 924 27808 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 29552 0 1 8976
box 29552 8976 29752 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 29552 0 1 924
box 29552 924 29752 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 31496 0 1 8976
box 31496 8976 31696 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 31496 0 1 924
box 31496 924 31696 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 33440 0 1 8976
box 33440 8976 33640 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 33440 0 1 924
box 33440 924 33640 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 35384 0 1 8976
box 35384 8976 35584 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 35384 0 1 924
box 35384 924 35584 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 37328 0 1 8976
box 37328 8976 37528 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 37328 0 1 924
box 37328 924 37528 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 39272 0 1 8976
box 39272 8976 39472 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 39272 0 1 924
box 39272 924 39472 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 41216 0 1 8976
box 41216 8976 41416 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 41216 0 1 924
box 41216 924 41416 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 43160 0 1 8976
box 43160 8976 43360 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 43160 0 1 924
box 43160 924 43360 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 45104 0 1 8976
box 45104 8976 45304 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 45104 0 1 924
box 45104 924 45304 1000
use RPLYBS_cut_M1M4_2x1 
transform 1 0 47048 0 1 8976
box 47048 8976 47248 9052
use RPLYBS_cut_M3M4_2x1 
transform 1 0 47048 0 1 924
box 47048 924 47248 1000
use RPLYBS_cut_M1M2_2x1 
transform 1 0 2344 0 1 12144
box 2344 12144 2528 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 2336 0 1 19076
box 2336 19076 2536 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 4288 0 1 12144
box 4288 12144 4472 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 4280 0 1 19076
box 4280 19076 4480 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 6232 0 1 12144
box 6232 12144 6416 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 6224 0 1 19076
box 6224 19076 6424 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 8176 0 1 12144
box 8176 12144 8360 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 8168 0 1 19076
box 8168 19076 8368 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 10120 0 1 12144
box 10120 12144 10304 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 10112 0 1 19076
box 10112 19076 10312 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 12064 0 1 12144
box 12064 12144 12248 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 12056 0 1 19076
box 12056 19076 12256 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 14008 0 1 12144
box 14008 12144 14192 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 14000 0 1 19076
box 14000 19076 14200 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 15952 0 1 12144
box 15952 12144 16136 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 15944 0 1 19076
box 15944 19076 16144 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 17896 0 1 12144
box 17896 12144 18080 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 17888 0 1 19076
box 17888 19076 18088 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 19840 0 1 12144
box 19840 12144 20024 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 19832 0 1 19076
box 19832 19076 20032 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 21784 0 1 12144
box 21784 12144 21968 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 21776 0 1 19076
box 21776 19076 21976 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 23728 0 1 12144
box 23728 12144 23912 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 23720 0 1 19076
box 23720 19076 23920 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 25672 0 1 12144
box 25672 12144 25856 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 25664 0 1 19076
box 25664 19076 25864 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 27616 0 1 12144
box 27616 12144 27800 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 27608 0 1 19076
box 27608 19076 27808 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 29560 0 1 12144
box 29560 12144 29744 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 29552 0 1 19076
box 29552 19076 29752 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 31504 0 1 12144
box 31504 12144 31688 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 31496 0 1 19076
box 31496 19076 31696 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 33448 0 1 12144
box 33448 12144 33632 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 33440 0 1 19076
box 33440 19076 33640 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 35392 0 1 12144
box 35392 12144 35576 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 35384 0 1 19076
box 35384 19076 35584 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 37336 0 1 12144
box 37336 12144 37520 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 37328 0 1 19076
box 37328 19076 37528 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 39280 0 1 12144
box 39280 12144 39464 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 39272 0 1 19076
box 39272 19076 39472 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 41224 0 1 12144
box 41224 12144 41408 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 41216 0 1 19076
box 41216 19076 41416 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 43168 0 1 12144
box 43168 12144 43352 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 43160 0 1 19076
box 43160 19076 43360 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 45112 0 1 12144
box 45112 12144 45296 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 45104 0 1 19076
box 45104 19076 45304 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 47056 0 1 12144
box 47056 12144 47240 12212
use RPLYBS_cut_M2M3_2x1 
transform 1 0 47048 0 1 19076
box 47048 19076 47248 19152
use RPLYBS_cut_M1M2_2x1 
transform 1 0 1392 0 1 11968
box 1392 11968 1576 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 1384 0 1 20104
box 1384 20104 1584 20180
use RPLYBS_cut_M1M2_2x1 
transform 1 0 3336 0 1 11968
box 3336 11968 3520 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 3328 0 1 20104
box 3328 20104 3528 20180
use RPLYBS_cut_M1M2_2x1 
transform 1 0 5280 0 1 11968
box 5280 11968 5464 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 5272 0 1 20104
box 5272 20104 5472 20180
use RPLYBS_cut_M1M2_2x1 
transform 1 0 7224 0 1 11968
box 7224 11968 7408 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 7216 0 1 20104
box 7216 20104 7416 20180
use RPLYBS_cut_M1M2_2x1 
transform 1 0 11112 0 1 11968
box 11112 11968 11296 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 11104 0 1 20104
box 11104 20104 11304 20180
use RPLYBS_cut_M1M2_2x1 
transform 1 0 13056 0 1 11968
box 13056 11968 13240 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 13048 0 1 20104
box 13048 20104 13248 20180
use RPLYBS_cut_M1M2_2x1 
transform 1 0 15000 0 1 11968
box 15000 11968 15184 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 14992 0 1 20104
box 14992 20104 15192 20180
use RPLYBS_cut_M1M2_2x1 
transform 1 0 16944 0 1 11968
box 16944 11968 17128 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 16936 0 1 20104
box 16936 20104 17136 20180
use RPLYBS_cut_M1M2_2x1 
transform 1 0 18888 0 1 11968
box 18888 11968 19072 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 18880 0 1 20104
box 18880 20104 19080 20180
use RPLYBS_cut_M1M2_2x1 
transform 1 0 20832 0 1 11968
box 20832 11968 21016 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 20824 0 1 20104
box 20824 20104 21024 20180
use RPLYBS_cut_M1M2_2x1 
transform 1 0 22776 0 1 11968
box 22776 11968 22960 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 22768 0 1 20104
box 22768 20104 22968 20180
use RPLYBS_cut_M1M2_2x1 
transform 1 0 24720 0 1 11968
box 24720 11968 24904 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 24712 0 1 20104
box 24712 20104 24912 20180
use RPLYBS_cut_M1M2_2x1 
transform 1 0 28608 0 1 11968
box 28608 11968 28792 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 28600 0 1 20104
box 28600 20104 28800 20180
use RPLYBS_cut_M1M2_2x1 
transform 1 0 30552 0 1 11968
box 30552 11968 30736 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 30544 0 1 20104
box 30544 20104 30744 20180
use RPLYBS_cut_M1M2_2x1 
transform 1 0 32496 0 1 11968
box 32496 11968 32680 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 32488 0 1 20104
box 32488 20104 32688 20180
use RPLYBS_cut_M1M2_2x1 
transform 1 0 34440 0 1 11968
box 34440 11968 34624 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 34432 0 1 20104
box 34432 20104 34632 20180
use RPLYBS_cut_M1M2_2x1 
transform 1 0 9168 0 1 11968
box 9168 11968 9352 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 9160 0 1 20544
box 9160 20544 9360 20620
use RPLYBS_cut_M1M2_2x1 
transform 1 0 26664 0 1 11968
box 26664 11968 26848 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 26656 0 1 20544
box 26656 20544 26856 20620
use RPLYBS_cut_M1M2_2x1 
transform 1 0 38328 0 1 11968
box 38328 11968 38512 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 38320 0 1 20768
box 38320 20768 38520 20844
use RPLYBS_cut_M1M2_2x1 
transform 1 0 40272 0 1 11968
box 40272 11968 40456 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 40264 0 1 20992
box 40264 20992 40464 21068
use RPLYBS_cut_M1M2_2x1 
transform 1 0 42216 0 1 11968
box 42216 11968 42400 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 42208 0 1 21216
box 42208 21216 42408 21292
use RPLYBS_cut_M1M2_2x1 
transform 1 0 44160 0 1 11968
box 44160 11968 44344 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 44152 0 1 21440
box 44152 21440 44352 21516
use RPLYBS_cut_M1M2_2x1 
transform 1 0 46104 0 1 11968
box 46104 11968 46288 12036
use RPLYBS_cut_M2M3_2x1 
transform 1 0 46096 0 1 21664
box 46096 21664 46296 21740
use RPLYBS_cut_M1M3_2x1 
transform 1 0 2328 0 1 2640
box 2328 2640 2528 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 4272 0 1 2640
box 4272 2640 4472 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 6216 0 1 2640
box 6216 2640 6416 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 8160 0 1 2640
box 8160 2640 8360 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 10104 0 1 2640
box 10104 2640 10304 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 12048 0 1 2640
box 12048 2640 12248 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 13992 0 1 2640
box 13992 2640 14192 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 15936 0 1 2640
box 15936 2640 16136 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 17880 0 1 2640
box 17880 2640 18080 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 19824 0 1 2640
box 19824 2640 20024 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 21768 0 1 2640
box 21768 2640 21968 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 23712 0 1 2640
box 23712 2640 23912 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 25656 0 1 2640
box 25656 2640 25856 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 27600 0 1 2640
box 27600 2640 27800 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 29544 0 1 2640
box 29544 2640 29744 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 31488 0 1 2640
box 31488 2640 31688 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 33432 0 1 2640
box 33432 2640 33632 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 35376 0 1 2640
box 35376 2640 35576 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 37320 0 1 2640
box 37320 2640 37520 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 39264 0 1 2640
box 39264 2640 39464 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 41208 0 1 2640
box 41208 2640 41408 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 43152 0 1 2640
box 43152 2640 43352 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 45096 0 1 2640
box 45096 2640 45296 2716
use RPLYBS_cut_M1M3_2x1 
transform 1 0 47040 0 1 2640
box 47040 2640 47240 2716
<< labels >>
flabel m2 s 0 924 46656 1076 0 FreeSans 400 0 0 0 VBP
port 1 nsew
flabel m2 s 0 19076 46656 19228 0 FreeSans 400 0 0 0 VCP
port 2 nsew
flabel locali s 47868 336 48168 19816 0 FreeSans 400 0 0 0 AVDD
port 11 nsew
flabel m2 s 1384 20104 34632 20256 0 FreeSans 400 0 0 0 IBP_A
port 3 nsew
flabel m2 s 9160 20544 26856 20696 0 FreeSans 400 0 0 0 IBP_B
port 4 nsew
flabel m2 s 38320 20768 38520 20920 0 FreeSans 400 0 0 0 IBP_1U<4>
port 6 nsew
flabel m2 s 40264 20992 40464 21144 0 FreeSans 400 0 0 0 IBP_1U<3>
port 7 nsew
flabel m2 s 42208 21216 42408 21368 0 FreeSans 400 0 0 0 IBP_1U<2>
port 8 nsew
flabel m2 s 44152 21440 44352 21592 0 FreeSans 400 0 0 0 IBP_1U<1>
port 9 nsew
flabel m2 s 46096 21664 46296 21816 0 FreeSans 400 0 0 0 IBP_1U<0>
port 10 nsew
flabel locali s 16 16 48488 128 0 FreeSans 400 0 0 0 VSS
port 12 nsew
flabel locali s 36384 11968 37104 12056 0 FreeSans 400 0 0 0 IBP_1U<5>
port 5 nsew
flabel m2 s 0 2640 216 2728 0 FreeSans 400 0 0 0 PWRUP_N
port 13 nsew
<< end >>
