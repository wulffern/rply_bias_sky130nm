
.subckt PCHCM D G S B
X1 D G S B PCH S=4
.ends

.subckt NCHCM D G S B
X1 D G S B NCH S=4
.ends

.subckt NCHA D G S B
X1 D G S B NCH M=2
.ends


.subckt PCHA D G S B
X1 D G S B PCH M=4
.ends


.subckt PCM OUT VCP VBP AVDD PWRUP_N
X1DMY0 AVDD AVDD AVDD AVDD PCH
X1SW SWD PWRUP_N AVDD AVDD PCHA
X1CM DCM VBP SWD AVDD PCHCM
X1CA OUT VCP DCM AVDD PCHA
X1DMY1 AVDD AVDD AVDD AVDD PCH
.ends

.subckt PMIRR VBP VCP IBP_A IBP_B  IBP_1U<5> IBP_1U<4> IBP_1U<3> IBP_1U<2> IBP_1U<1> IBP_1U<0> AVDD VSS PWRUP_N
XA01 IBP_A VCP VBP AVDD PWRUP_N PCM M=4
XB02 IBP_B VCP VBP AVDD PWRUP_N PCM M=1
XC03 IBP_A VCP VBP AVDD PWRUP_N PCM M=4
XD04 IBP_A VCP VBP AVDD PWRUP_N PCM M=4
XB02a IBP_B VCP VBP AVDD PWRUP_N PCM M=1
XF06 IBP_A VCP VBP AVDD PWRUP_N PCM M=4
XG05a VBP VCP VBP AVDD PWRUP_N PCM
XG05 IBP_1U<5> VCP VBP AVDD PWRUP_N PCM
XG07 IBP_1U<4> VCP VBP AVDD PWRUP_N PCM
XH08 IBP_1U<3> VCP VBP AVDD PWRUP_N PCM
XI09 IBP_1U<2> VCP VBP AVDD PWRUP_N PCM
XJ10 IBP_1U<1> VCP VBP AVDD PWRUP_N PCM
XK11 IBP_1U<0> VCP VBP AVDD PWRUP_N PCM
.ends
