magic
tech sky130B
magscale 1 2
timestamp 1675206000
<< checkpaint >>
rect 0 0 1944 792
<< pdiff >>
rect 468 132 1188 220
rect 468 220 1188 308
rect 468 308 1188 396
rect 468 396 1188 484
rect 468 484 1188 572
rect 468 572 1188 660
<< ntap >>
rect -108 -44 108 44
rect 1836 -44 2052 44
rect -108 44 108 132
rect 1836 44 2052 132
rect -108 132 108 220
rect 1836 132 2052 220
rect -108 220 108 308
rect 1836 220 2052 308
rect -108 308 108 396
rect 1836 308 2052 396
rect -108 396 108 484
rect 1836 396 2052 484
rect -108 484 108 572
rect 1836 484 2052 572
rect -108 572 108 660
rect 1836 572 2052 660
rect -108 660 108 748
rect 1836 660 2052 748
rect -108 748 108 836
rect 1836 748 2052 836
<< poly >>
rect 396 -36 1620 36
rect 396 228 1620 300
rect 396 492 1620 564
rect 396 756 1620 828
rect 1404 220 1620 308
rect 1404 484 1620 572
<< locali >>
rect 1404 484 1620 572
rect -108 -44 108 44
rect 1836 -44 2052 44
rect -108 44 108 132
rect 1836 44 2052 132
rect -108 132 108 220
rect 324 132 1188 220
rect 324 132 1188 220
rect 1836 132 2052 220
rect -108 220 108 308
rect 1836 484 2052 572
rect 324 220 396 308
rect 1404 220 1620 308
rect 1836 220 2052 308
rect -108 308 108 396
rect 324 308 396 396
rect 468 308 1188 396
rect 468 308 1188 396
rect 1476 308 1548 396
rect 1836 308 2052 396
rect -108 396 108 484
rect 324 396 396 484
rect 468 396 1188 484
rect 1476 396 1548 484
rect 1836 396 2052 484
rect -108 484 108 572
rect 324 484 396 572
rect 1404 484 1620 572
rect 1836 484 2052 572
rect -108 572 108 660
rect 324 572 1188 660
rect 1836 572 2052 660
rect -108 660 108 748
rect 1836 660 2052 748
rect -108 748 108 836
rect 1836 748 2052 836
<< pcontact >>
rect 1428 242 1476 264
rect 1428 264 1476 286
rect 1476 242 1548 264
rect 1476 264 1548 286
rect 1548 242 1596 264
rect 1548 264 1596 286
rect 1428 506 1476 528
rect 1428 528 1476 550
rect 1476 506 1548 528
rect 1476 528 1548 550
rect 1548 506 1596 528
rect 1548 528 1596 550
<< ntapc >>
rect -36 132 36 220
rect 1908 132 1980 220
rect -36 220 36 308
rect 1908 220 1980 308
rect -36 308 36 396
rect 1908 308 1980 396
rect -36 396 36 484
rect 1908 396 1980 484
rect -36 484 36 572
rect 1908 484 1980 572
rect -36 572 36 660
rect 1908 572 1980 660
<< pdcontact >>
rect 492 154 540 176
rect 492 176 540 198
rect 540 154 612 176
rect 540 176 612 198
rect 612 154 684 176
rect 612 176 684 198
rect 684 154 756 176
rect 684 176 756 198
rect 756 154 828 176
rect 756 176 828 198
rect 828 154 900 176
rect 828 176 900 198
rect 900 154 972 176
rect 900 176 972 198
rect 972 154 1044 176
rect 972 176 1044 198
rect 1044 154 1116 176
rect 1044 176 1116 198
rect 1116 154 1164 176
rect 1116 176 1164 198
rect 492 330 540 352
rect 492 352 540 374
rect 540 330 612 352
rect 540 352 612 374
rect 612 330 684 352
rect 612 352 684 374
rect 684 330 756 352
rect 684 352 756 374
rect 756 330 828 352
rect 756 352 828 374
rect 828 330 900 352
rect 828 352 900 374
rect 900 330 972 352
rect 900 352 972 374
rect 972 330 1044 352
rect 972 352 1044 374
rect 1044 330 1116 352
rect 1044 352 1116 374
rect 1116 330 1164 352
rect 1116 352 1164 374
rect 492 418 540 440
rect 492 440 540 462
rect 540 418 612 440
rect 540 440 612 462
rect 612 418 684 440
rect 612 440 684 462
rect 684 418 756 440
rect 684 440 756 462
rect 756 418 828 440
rect 756 440 828 462
rect 828 418 900 440
rect 828 440 900 462
rect 900 418 972 440
rect 900 440 972 462
rect 972 418 1044 440
rect 972 440 1044 462
rect 1044 418 1116 440
rect 1044 440 1116 462
rect 1116 418 1164 440
rect 1116 440 1164 462
rect 492 594 540 616
rect 492 616 540 638
rect 540 594 612 616
rect 540 616 612 638
rect 612 594 684 616
rect 612 616 684 638
rect 684 594 756 616
rect 684 616 756 638
rect 756 594 828 616
rect 756 616 828 638
rect 828 594 900 616
rect 828 616 900 638
rect 900 594 972 616
rect 900 616 972 638
rect 972 594 1044 616
rect 972 616 1044 638
rect 1044 594 1116 616
rect 1044 616 1116 638
rect 1116 594 1164 616
rect 1116 616 1164 638
<< nwell >>
rect -180 -132 2124 924
<< labels >>
flabel locali s 1404 484 1620 572 0 FreeSans 400 0 0 0 G
port 2 nsew
flabel locali s 324 132 1188 220 0 FreeSans 400 0 0 0 S
port 3 nsew
flabel locali s 1836 484 2052 572 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel locali s 468 308 1188 396 0 FreeSans 400 0 0 0 D
port 1 nsew
<< end >>
