
*-------------------------------------------------------------
* RPLYBS_PCH <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT RPLYBS_PCH D G S B
XMM1 D G S B sky130_fd_pr__pfet_01v8  l=0.36  nf=2  w=3.6*nf  
.ENDS

*-------------------------------------------------------------
* RPLYBS_NCH <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT RPLYBS_NCH D G S B
XMM1 D G S B sky130_fd_pr__nfet_01v8  l=0.36  nf=2  w=3.6*nf  
.ENDS

*-------------------------------------------------------------
* RPLYBS_PCHCM <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT RPLYBS_PCHCM D G S B
X1_S0 D_S0 G S B RPLYBS_PCH
X1_S1 D_S1 G D_S0 B RPLYBS_PCH
X1_S2 D_S2 G D_S1 B RPLYBS_PCH
X1_S3 D G D_S2 B RPLYBS_PCH
.ENDS

*-------------------------------------------------------------
* RPLYBS_NCHCM <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT RPLYBS_NCHCM D G S B
X1_S0 D_S0 G S B RPLYBS_NCH
X1_S1 D_S1 G D_S0 B RPLYBS_NCH
X1_S2 D_S2 G D_S1 B RPLYBS_NCH
X1_S3 D G D_S2 B RPLYBS_NCH
.ENDS

*-------------------------------------------------------------
* RPLYBS_PCHA <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT RPLYBS_PCHA D G S B
X10 D G S B RPLYBS_PCH
X11 D G S B RPLYBS_PCH
X12 D G S B RPLYBS_PCH
X13 D G S B RPLYBS_PCH
.ENDS

*-------------------------------------------------------------
* RPLYBS_NCHA <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT RPLYBS_NCHA D G S B
X10 D G S B RPLYBS_NCH
X11 D G S B RPLYBS_NCH
.ENDS

*-------------------------------------------------------------
* RPLYBS_PCM <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT RPLYBS_PCM OUT VCP VBP AVDD PWRUP_N
X1DMY0 AVDD AVDD AVDD AVDD RPLYBS_PCH
X1SW SWD PWRUP_N AVDD AVDD RPLYBS_PCHA
X1CM DCM VBP SWD AVDD RPLYBS_PCHCM
X1CA OUT VCP DCM AVDD RPLYBS_PCHA
X1DMY1 AVDD AVDD AVDD AVDD RPLYBS_PCH
.ENDS

*-------------------------------------------------------------
* RPLYBS_PMIRR <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT RPLYBS_PMIRR VBP VCP IBP_A IBP_B IBP_1U_5 IBP_1U_4 IBP_1U_3 IBP_1U_2 IBP_1U_1 IBP_1U_0 AVDD VSS PWRUP_N
XA010 IBP_A VCP VBP AVDD PWRUP_N RPLYBS_PCM
XA011 IBP_A VCP VBP AVDD PWRUP_N RPLYBS_PCM
XA012 IBP_A VCP VBP AVDD PWRUP_N RPLYBS_PCM
XA013 IBP_A VCP VBP AVDD PWRUP_N RPLYBS_PCM
XB020 IBP_B VCP VBP AVDD PWRUP_N RPLYBS_PCM
XC030 IBP_A VCP VBP AVDD PWRUP_N RPLYBS_PCM
XC031 IBP_A VCP VBP AVDD PWRUP_N RPLYBS_PCM
XC032 IBP_A VCP VBP AVDD PWRUP_N RPLYBS_PCM
XC033 IBP_A VCP VBP AVDD PWRUP_N RPLYBS_PCM
XD040 IBP_A VCP VBP AVDD PWRUP_N RPLYBS_PCM
XD041 IBP_A VCP VBP AVDD PWRUP_N RPLYBS_PCM
XD042 IBP_A VCP VBP AVDD PWRUP_N RPLYBS_PCM
XD043 IBP_A VCP VBP AVDD PWRUP_N RPLYBS_PCM
XB02a0 IBP_B VCP VBP AVDD PWRUP_N RPLYBS_PCM
XF060 IBP_A VCP VBP AVDD PWRUP_N RPLYBS_PCM
XF061 IBP_A VCP VBP AVDD PWRUP_N RPLYBS_PCM
XF062 IBP_A VCP VBP AVDD PWRUP_N RPLYBS_PCM
XF063 IBP_A VCP VBP AVDD PWRUP_N RPLYBS_PCM
XG05a VBP VCP VBP AVDD PWRUP_N RPLYBS_PCM
XG05 IBP_1U_5 VCP VBP AVDD PWRUP_N RPLYBS_PCM
XG07 IBP_1U_4 VCP VBP AVDD PWRUP_N RPLYBS_PCM
XH08 IBP_1U_3 VCP VBP AVDD PWRUP_N RPLYBS_PCM
XI09 IBP_1U_2 VCP VBP AVDD PWRUP_N RPLYBS_PCM
XJ10 IBP_1U_1 VCP VBP AVDD PWRUP_N RPLYBS_PCM
XK11 IBP_1U_0 VCP VBP AVDD PWRUP_N RPLYBS_PCM
.ENDS
