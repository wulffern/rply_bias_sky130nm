magic
tech sky130B
magscale 1 2
timestamp 1675206000
<< checkpaint >>
rect 0 0 1944 1584
<< locali >>
rect 828 308 1248 368
rect 828 1100 1248 1160
rect 1248 308 1308 1160
rect 1482 484 1542 1364
rect 324 132 756 192
rect 324 924 756 984
rect 324 132 384 984
rect -108 220 108 308
rect 468 308 1188 396
rect 1404 484 1620 572
rect 324 132 1188 220
use RPLYBS_NCH X10
transform 1 0 0 0 1 0
box 0 0 1944 792
use RPLYBS_NCH X11
transform 1 0 0 0 1 792
box 0 792 1944 1584
<< labels >>
flabel locali s -108 220 108 308 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel locali s 468 308 1188 396 0 FreeSans 400 0 0 0 D
port 1 nsew
flabel locali s 1404 484 1620 572 0 FreeSans 400 0 0 0 G
port 2 nsew
flabel locali s 324 132 1188 220 0 FreeSans 400 0 0 0 S
port 3 nsew
<< end >>
