magic
tech sky130B
magscale 1 2
timestamp 1672527600
<< checkpaint >>
rect 0 0 1944 6336
<< locali >>
rect 756 924 1248 984
rect 828 308 1248 368
rect 1248 308 1308 984
rect 756 1716 1248 1776
rect 828 1100 1248 1160
rect 1248 1100 1308 1776
rect 756 2508 1248 2568
rect 828 1892 1248 1952
rect 1248 1892 1308 2568
rect 756 3300 1248 3360
rect 828 2684 1248 2744
rect 1248 2684 1308 3360
rect 756 4092 1248 4152
rect 828 3476 1248 3536
rect 1248 3476 1308 4152
rect 756 4884 1248 4944
rect 828 4268 1248 4328
rect 1248 4268 1308 4944
rect 756 5676 1248 5736
rect 828 5060 1248 5120
rect 1248 5060 1308 5736
rect 828 5852 1248 5912
rect 1248 5852 1308 5912
rect 1482 484 1542 6116
rect -108 220 108 308
rect 468 5852 1188 5940
rect 1404 484 1620 572
rect 324 132 1188 220
use RPLYBS_NCH X1_S0
transform 1 0 0 0 1 0
box 0 0 1944 792
use RPLYBS_NCH X1_S1
transform 1 0 0 0 1 792
box 0 792 1944 1584
use RPLYBS_NCH X1_S2
transform 1 0 0 0 1 1584
box 0 1584 1944 2376
use RPLYBS_NCH X1_S3
transform 1 0 0 0 1 2376
box 0 2376 1944 3168
use RPLYBS_NCH X1_S4
transform 1 0 0 0 1 3168
box 0 3168 1944 3960
use RPLYBS_NCH X1_S5
transform 1 0 0 0 1 3960
box 0 3960 1944 4752
use RPLYBS_NCH X1_S6
transform 1 0 0 0 1 4752
box 0 4752 1944 5544
use RPLYBS_NCH X1_S7
transform 1 0 0 0 1 5544
box 0 5544 1944 6336
<< labels >>
flabel locali s -108 220 108 308 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel locali s 468 5852 1188 5940 0 FreeSans 400 0 0 0 D
port 1 nsew
flabel locali s 1404 484 1620 572 0 FreeSans 400 0 0 0 G
port 2 nsew
flabel locali s 324 132 1188 220 0 FreeSans 400 0 0 0 S
port 3 nsew
<< end >>
