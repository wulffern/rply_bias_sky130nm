*RPLY_BIAS_SKY130A/RPLY_BIAS
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/RPLY_BIAS_lpe.spi
#else
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_CAP_10_lpe.spi
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_CAP_20_lpe.spi
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_PCHDLCM_lpe.spi
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_PCHL_lpe.spi
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_PCHDL_lpe.spi
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_NCHDLCM_lpe.spi
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_NCHDL_lpe.spi
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_PCHDLA_lpe.spi
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_NCHL_lpe.spi
.include ../../../work/xsch/RPLY_BIAS.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
#ifdef Debug
.option reltol=1e-3 srcsteps=1 ramptime=10n noopiter keepopinfo gmin=1e-12 method=gear
#else
.option reltol=1e-6 srcsteps=1 ramptime=10n noopiter gmin=1e-15
#endif

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

.param T_END = {1u}
.csparam T_END = {T_END}+100p

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  0  dc  {AVDD}
VPWR  PWRUP_1V8  0 dc {AVDD}

VLST LPI LPO dc 0


*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VDD_1V8 VSS PWRUP_1V8 LPI LPO
+ IBP_1U<3>,IBP_1U<2>,IBP_1U<1>,IBP_1U<0> T_OP T_ON RPLY_BIAS

*-----------------------------------------------------------------
* STASH
*-----------------------------------------------------------------

V3 IBP_1U<3> 0 dc {AVDD/2}
V2 IBP_1U<2> 0 dc {AVDD/2}
V1 IBP_1U<1> 0 dc {AVDD/2}
V0 IBP_1U<0> 0 dc {AVDD/2}

* Save temperature to transient
B5 temp 0 v=temper
*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
*.save all
#else
.save v(VDD_1V8) v(VSS) v(PWRUP_1V8) v(LPI) v(LPO) v(IBP_1U) i(v1)
+ v(XDUT.VD1) v(XDUT.VD2) v(XDUT.VR1) v(D_VD) v(D_VD_REF) v(D_VD_ERR)
+ v(V_OFF) i(VDD)
+ v(xdut.xota.vs1)
+ v(xdut.xota.vbp2)
+ v(xdut.xota.vo_ls)
+ v(xdut.ibp_2u)
+ v(xdut.xota.vs)
+ v(xdut.xota.vbp1)
+ v(xdut.xota.vbp2)
+ v(xdut.xota.vbp3)
+ v(xdut.xota.vbn1)
+ v(xdut.xota.vbn2)
+ v(xdut.vip)
+ v(xdut.vin)
+ v(xdut.xota.vstart)
+ v(xdut.xota.vstarted)
*+ v(xdut.xota.vin_ls) v(xdut.xota.vip_ls) v(xdut.xota.vs) v(xdut.xota.vbpb) v(xdut.xota.vbp)
+ v(t_op) v(t_on)
+ v(temp)
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set ng_nomodcheck
set keepopinfo
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 10n 1u 0


dc TEMP -40 125 5

write
#ifdef Debug


*quit
#else

quit
#endif
.endc
